module bitmap_rom (
    input wire [6:0] x,
    input wire [6:0] y,
    output wire [2:0] pixel
);

  reg [2:0] mem[2047:0];
  initial begin
    mem[0] = 3'd0;
    mem[1] = 3'd0;
    mem[2] = 3'd0;
    mem[3] = 3'd0;
    mem[4] = 3'd0;
    mem[5] = 3'd0;
    mem[6] = 3'd0;
    mem[7] = 3'd0;
    mem[8] = 3'd0;
    mem[9] = 3'd0;
    mem[10] = 3'd0;
    mem[11] = 3'd0;
    mem[12] = 3'd0;
    mem[13] = 3'd0;
    mem[14] = 3'd0;
    mem[15] = 3'd0;
    mem[16] = 3'd0;
    mem[17] = 3'd0;
    mem[18] = 3'd0;
    mem[19] = 3'd0;
    mem[20] = 3'd0;
    mem[21] = 3'd0;
    mem[22] = 3'd7;
    mem[23] = 3'd7;
    mem[24] = 3'd7;
    mem[25] = 3'd0;
    mem[26] = 3'd0;
    mem[27] = 3'd0;
    mem[28] = 3'd0;
    mem[29] = 3'd0;
    mem[30] = 3'd0;
    mem[31] = 3'd0;
    mem[32] = 3'd0;
    mem[33] = 3'd0;
    mem[34] = 3'd0;
    mem[35] = 3'd0;
    mem[36] = 3'd0;
    mem[37] = 3'd0;
    mem[38] = 3'd7;
    mem[39] = 3'd7;
    mem[40] = 3'd7;
    mem[41] = 3'd0;
    mem[42] = 3'd0;
    mem[43] = 3'd0;
    mem[44] = 3'd0;
    mem[45] = 3'd0;
    mem[46] = 3'd0;
    mem[47] = 3'd0;
    mem[48] = 3'd0;
    mem[49] = 3'd0;
    mem[50] = 3'd0;
    mem[51] = 3'd0;
    mem[52] = 3'd0;
    mem[53] = 3'd7;
    mem[54] = 3'd7;
    mem[55] = 3'd7;
    mem[56] = 3'd7;
    mem[57] = 3'd7;
    mem[58] = 3'd0;
    mem[59] = 3'd0;
    mem[60] = 3'd0;
    mem[61] = 3'd0;
    mem[62] = 3'd0;
    mem[63] = 3'd0;
    mem[64] = 3'd0;
    mem[65] = 3'd0;
    mem[66] = 3'd0;
    mem[67] = 3'd0;
    mem[68] = 3'd0;
    mem[69] = 3'd7;
    mem[70] = 3'd7;
    mem[71] = 3'd7;
    mem[72] = 3'd7;
    mem[73] = 3'd7;
    mem[74] = 3'd0;
    mem[75] = 3'd0;
    mem[76] = 3'd0;
    mem[77] = 3'd0;
    mem[78] = 3'd0;
    mem[79] = 3'd0;
    mem[80] = 3'd0;
    mem[81] = 3'd0;
    mem[82] = 3'd0;
    mem[83] = 3'd0;
    mem[84] = 3'd0;
    mem[85] = 3'd7;
    mem[86] = 3'd7;
    mem[87] = 3'd7;
    mem[88] = 3'd7;
    mem[89] = 3'd7;
    mem[90] = 3'd7;
    mem[91] = 3'd0;
    mem[92] = 3'd0;
    mem[93] = 3'd0;
    mem[94] = 3'd0;
    mem[95] = 3'd0;
    mem[96] = 3'd0;
    mem[97] = 3'd0;
    mem[98] = 3'd0;
    mem[99] = 3'd0;
    mem[100] = 3'd7;
    mem[101] = 3'd7;
    mem[102] = 3'd7;
    mem[103] = 3'd7;
    mem[104] = 3'd7;
    mem[105] = 3'd7;
    mem[106] = 3'd7;
    mem[107] = 3'd0;
    mem[108] = 3'd0;
    mem[109] = 3'd0;
    mem[110] = 3'd0;
    mem[111] = 3'd0;
    mem[112] = 3'd0;
    mem[113] = 3'd0;
    mem[114] = 3'd0;
    mem[115] = 3'd0;
    mem[116] = 3'd7;
    mem[117] = 3'd7;
    mem[118] = 3'd7;
    mem[119] = 3'd7;
    mem[120] = 3'd7;
    mem[121] = 3'd7;
    mem[122] = 3'd7;
    mem[123] = 3'd0;
    mem[124] = 3'd0;
    mem[125] = 3'd0;
    mem[126] = 3'd0;
    mem[127] = 3'd0;
    mem[128] = 3'd0;
    mem[129] = 3'd0;
    mem[130] = 3'd0;
    mem[131] = 3'd0;
    mem[132] = 3'd7;
    mem[133] = 3'd7;
    mem[134] = 3'd7;
    mem[135] = 3'd7;
    mem[136] = 3'd7;
    mem[137] = 3'd7;
    mem[138] = 3'd7;
    mem[139] = 3'd0;
    mem[140] = 3'd0;
    mem[141] = 3'd0;
    mem[142] = 3'd0;
    mem[143] = 3'd0;
    mem[144] = 3'd0;
    mem[145] = 3'd0;
    mem[146] = 3'd0;
    mem[147] = 3'd0;
    mem[148] = 3'd7;
    mem[149] = 3'd7;
    mem[150] = 3'd7;
    mem[151] = 3'd7;
    mem[152] = 3'd7;
    mem[153] = 3'd7;
    mem[154] = 3'd7;
    mem[155] = 3'd7;
    mem[156] = 3'd0;
    mem[157] = 3'd0;
    mem[158] = 3'd0;
    mem[159] = 3'd0;
    mem[160] = 3'd0;
    mem[161] = 3'd0;
    mem[162] = 3'd0;
    mem[163] = 3'd7;
    mem[164] = 3'd7;
    mem[165] = 3'd7;
    mem[166] = 3'd7;
    mem[167] = 3'd7;
    mem[168] = 3'd7;
    mem[169] = 3'd7;
    mem[170] = 3'd7;
    mem[171] = 3'd7;
    mem[172] = 3'd0;
    mem[173] = 3'd0;
    mem[174] = 3'd0;
    mem[175] = 3'd0;
    mem[176] = 3'd0;
    mem[177] = 3'd0;
    mem[178] = 3'd0;
    mem[179] = 3'd7;
    mem[180] = 3'd7;
    mem[181] = 3'd7;
    mem[182] = 3'd7;
    mem[183] = 3'd7;
    mem[184] = 3'd7;
    mem[185] = 3'd7;
    mem[186] = 3'd7;
    mem[187] = 3'd7;
    mem[188] = 3'd0;
    mem[189] = 3'd0;
    mem[190] = 3'd0;
    mem[191] = 3'd0;
    mem[192] = 3'd0;
    mem[193] = 3'd0;
    mem[194] = 3'd0;
    mem[195] = 3'd7;
    mem[196] = 3'd7;
    mem[197] = 3'd7;
    mem[198] = 3'd0;
    mem[199] = 3'd0;
    mem[200] = 3'd0;
    mem[201] = 3'd7;
    mem[202] = 3'd7;
    mem[203] = 3'd7;
    mem[204] = 3'd0;
    mem[205] = 3'd0;
    mem[206] = 3'd0;
    mem[207] = 3'd0;
    mem[208] = 3'd0;
    mem[209] = 3'd0;
    mem[210] = 3'd0;
    mem[211] = 3'd7;
    mem[212] = 3'd7;
    mem[213] = 3'd7;
    mem[214] = 3'd0;
    mem[215] = 3'd0;
    mem[216] = 3'd0;
    mem[217] = 3'd7;
    mem[218] = 3'd7;
    mem[219] = 3'd7;
    mem[220] = 3'd0;
    mem[221] = 3'd0;
    mem[222] = 3'd0;
    mem[223] = 3'd0;
    mem[224] = 3'd0;
    mem[225] = 3'd0;
    mem[226] = 3'd0;
    mem[227] = 3'd7;
    mem[228] = 3'd7;
    mem[229] = 3'd7;
    mem[230] = 3'd0;
    mem[231] = 3'd0;
    mem[232] = 3'd0;
    mem[233] = 3'd0;
    mem[234] = 3'd7;
    mem[235] = 3'd7;
    mem[236] = 3'd7;
    mem[237] = 3'd0;
    mem[238] = 3'd0;
    mem[239] = 3'd0;
    mem[240] = 3'd0;
    mem[241] = 3'd0;
    mem[242] = 3'd7;
    mem[243] = 3'd7;
    mem[244] = 3'd7;
    mem[245] = 3'd0;
    mem[246] = 3'd0;
    mem[247] = 3'd0;
    mem[248] = 3'd0;
    mem[249] = 3'd0;
    mem[250] = 3'd7;
    mem[251] = 3'd7;
    mem[252] = 3'd7;
    mem[253] = 3'd0;
    mem[254] = 3'd0;
    mem[255] = 3'd0;
    mem[256] = 3'd0;
    mem[257] = 3'd0;
    mem[258] = 3'd7;
    mem[259] = 3'd7;
    mem[260] = 3'd7;
    mem[261] = 3'd0;
    mem[262] = 3'd0;
    mem[263] = 3'd0;
    mem[264] = 3'd0;
    mem[265] = 3'd0;
    mem[266] = 3'd7;
    mem[267] = 3'd7;
    mem[268] = 3'd7;
    mem[269] = 3'd0;
    mem[270] = 3'd0;
    mem[271] = 3'd0;
    mem[272] = 3'd0;
    mem[273] = 3'd0;
    mem[274] = 3'd7;
    mem[275] = 3'd7;
    mem[276] = 3'd7;
    mem[277] = 3'd0;
    mem[278] = 3'd0;
    mem[279] = 3'd0;
    mem[280] = 3'd0;
    mem[281] = 3'd0;
    mem[282] = 3'd0;
    mem[283] = 3'd7;
    mem[284] = 3'd7;
    mem[285] = 3'd0;
    mem[286] = 3'd0;
    mem[287] = 3'd0;
    mem[288] = 3'd0;
    mem[289] = 3'd0;
    mem[290] = 3'd7;
    mem[291] = 3'd7;
    mem[292] = 3'd0;
    mem[293] = 3'd0;
    mem[294] = 3'd0;
    mem[295] = 3'd0;
    mem[296] = 3'd0;
    mem[297] = 3'd0;
    mem[298] = 3'd0;
    mem[299] = 3'd7;
    mem[300] = 3'd7;
    mem[301] = 3'd0;
    mem[302] = 3'd0;
    mem[303] = 3'd0;
    mem[304] = 3'd0;
    mem[305] = 3'd0;
    mem[306] = 3'd7;
    mem[307] = 3'd7;
    mem[308] = 3'd0;
    mem[309] = 3'd0;
    mem[310] = 3'd0;
    mem[311] = 3'd0;
    mem[312] = 3'd0;
    mem[313] = 3'd0;
    mem[314] = 3'd0;
    mem[315] = 3'd7;
    mem[316] = 3'd7;
    mem[317] = 3'd0;
    mem[318] = 3'd0;
    mem[319] = 3'd0;
    mem[320] = 3'd0;
    mem[321] = 3'd0;
    mem[322] = 3'd7;
    mem[323] = 3'd7;
    mem[324] = 3'd0;
    mem[325] = 3'd0;
    mem[326] = 3'd0;
    mem[327] = 3'd0;
    mem[328] = 3'd0;
    mem[329] = 3'd0;
    mem[330] = 3'd0;
    mem[331] = 3'd7;
    mem[332] = 3'd7;
    mem[333] = 3'd0;
    mem[334] = 3'd0;
    mem[335] = 3'd0;
    mem[336] = 3'd0;
    mem[337] = 3'd0;
    mem[338] = 3'd7;
    mem[339] = 3'd7;
    mem[340] = 3'd0;
    mem[341] = 3'd0;
    mem[342] = 3'd0;
    mem[343] = 3'd0;
    mem[344] = 3'd0;
    mem[345] = 3'd0;
    mem[346] = 3'd0;
    mem[347] = 3'd7;
    mem[348] = 3'd7;
    mem[349] = 3'd7;
    mem[350] = 3'd0;
    mem[351] = 3'd0;
    mem[352] = 3'd0;
    mem[353] = 3'd0;
    mem[354] = 3'd7;
    mem[355] = 3'd7;
    mem[356] = 3'd0;
    mem[357] = 3'd0;
    mem[358] = 3'd0;
    mem[359] = 3'd0;
    mem[360] = 3'd0;
    mem[361] = 3'd0;
    mem[362] = 3'd0;
    mem[363] = 3'd0;
    mem[364] = 3'd7;
    mem[365] = 3'd7;
    mem[366] = 3'd0;
    mem[367] = 3'd0;
    mem[368] = 3'd0;
    mem[369] = 3'd7;
    mem[370] = 3'd7;
    mem[371] = 3'd7;
    mem[372] = 3'd0;
    mem[373] = 3'd0;
    mem[374] = 3'd0;
    mem[375] = 3'd0;
    mem[376] = 3'd0;
    mem[377] = 3'd0;
    mem[378] = 3'd0;
    mem[379] = 3'd0;
    mem[380] = 3'd7;
    mem[381] = 3'd7;
    mem[382] = 3'd0;
    mem[383] = 3'd0;
    mem[384] = 3'd0;
    mem[385] = 3'd7;
    mem[386] = 3'd7;
    mem[387] = 3'd0;
    mem[388] = 3'd0;
    mem[389] = 3'd0;
    mem[390] = 3'd0;
    mem[391] = 3'd0;
    mem[392] = 3'd0;
    mem[393] = 3'd0;
    mem[394] = 3'd0;
    mem[395] = 3'd0;
    mem[396] = 3'd7;
    mem[397] = 3'd7;
    mem[398] = 3'd0;
    mem[399] = 3'd0;
    mem[400] = 3'd0;
    mem[401] = 3'd7;
    mem[402] = 3'd7;
    mem[403] = 3'd0;
    mem[404] = 3'd0;
    mem[405] = 3'd0;
    mem[406] = 3'd0;
    mem[407] = 3'd0;
    mem[408] = 3'd0;
    mem[409] = 3'd0;
    mem[410] = 3'd0;
    mem[411] = 3'd0;
    mem[412] = 3'd7;
    mem[413] = 3'd7;
    mem[414] = 3'd0;
    mem[415] = 3'd0;
    mem[416] = 3'd0;
    mem[417] = 3'd7;
    mem[418] = 3'd7;
    mem[419] = 3'd0;
    mem[420] = 3'd0;
    mem[421] = 3'd0;
    mem[422] = 3'd0;
    mem[423] = 3'd0;
    mem[424] = 3'd0;
    mem[425] = 3'd0;
    mem[426] = 3'd0;
    mem[427] = 3'd0;
    mem[428] = 3'd7;
    mem[429] = 3'd7;
    mem[430] = 3'd0;
    mem[431] = 3'd0;
    mem[432] = 3'd0;
    mem[433] = 3'd7;
    mem[434] = 3'd7;
    mem[435] = 3'd7;
    mem[436] = 3'd7;
    mem[437] = 3'd7;
    mem[438] = 3'd7;
    mem[439] = 3'd7;
    mem[440] = 3'd7;
    mem[441] = 3'd0;
    mem[442] = 3'd0;
    mem[443] = 3'd0;
    mem[444] = 3'd7;
    mem[445] = 3'd7;
    mem[446] = 3'd0;
    mem[447] = 3'd0;
    mem[448] = 3'd0;
    mem[449] = 3'd7;
    mem[450] = 3'd7;
    mem[451] = 3'd7;
    mem[452] = 3'd7;
    mem[453] = 3'd7;
    mem[454] = 3'd7;
    mem[455] = 3'd7;
    mem[456] = 3'd7;
    mem[457] = 3'd0;
    mem[458] = 3'd0;
    mem[459] = 3'd0;
    mem[460] = 3'd7;
    mem[461] = 3'd7;
    mem[462] = 3'd0;
    mem[463] = 3'd0;
    mem[464] = 3'd0;
    mem[465] = 3'd7;
    mem[466] = 3'd7;
    mem[467] = 3'd7;
    mem[468] = 3'd7;
    mem[469] = 3'd7;
    mem[470] = 3'd7;
    mem[471] = 3'd7;
    mem[472] = 3'd7;
    mem[473] = 3'd0;
    mem[474] = 3'd0;
    mem[475] = 3'd0;
    mem[476] = 3'd7;
    mem[477] = 3'd7;
    mem[478] = 3'd0;
    mem[479] = 3'd0;
    mem[480] = 3'd0;
    mem[481] = 3'd7;
    mem[482] = 3'd7;
    mem[483] = 3'd7;
    mem[484] = 3'd7;
    mem[485] = 3'd7;
    mem[486] = 3'd7;
    mem[487] = 3'd7;
    mem[488] = 3'd7;
    mem[489] = 3'd0;
    mem[490] = 3'd0;
    mem[491] = 3'd0;
    mem[492] = 3'd0;
    mem[493] = 3'd7;
    mem[494] = 3'd0;
    mem[495] = 3'd0;
    mem[496] = 3'd0;
    mem[497] = 3'd7;
    mem[498] = 3'd7;
    mem[499] = 3'd7;
    mem[500] = 3'd7;
    mem[501] = 3'd7;
    mem[502] = 3'd7;
    mem[503] = 3'd7;
    mem[504] = 3'd7;
    mem[505] = 3'd0;
    mem[506] = 3'd0;
    mem[507] = 3'd0;
    mem[508] = 3'd0;
    mem[509] = 3'd7;
    mem[510] = 3'd0;
    mem[511] = 3'd0;
    mem[512] = 3'd0;
    mem[513] = 3'd7;
    mem[514] = 3'd7;
    mem[515] = 3'd7;
    mem[516] = 3'd7;
    mem[517] = 3'd7;
    mem[518] = 3'd7;
    mem[519] = 3'd7;
    mem[520] = 3'd7;
    mem[521] = 3'd0;
    mem[522] = 3'd0;
    mem[523] = 3'd0;
    mem[524] = 3'd0;
    mem[525] = 3'd7;
    mem[526] = 3'd7;
    mem[527] = 3'd0;
    mem[528] = 3'd0;
    mem[529] = 3'd7;
    mem[530] = 3'd7;
    mem[531] = 3'd7;
    mem[532] = 3'd7;
    mem[533] = 3'd7;
    mem[534] = 3'd7;
    mem[535] = 3'd7;
    mem[536] = 3'd7;
    mem[537] = 3'd0;
    mem[538] = 3'd0;
    mem[539] = 3'd0;
    mem[540] = 3'd0;
    mem[541] = 3'd7;
    mem[542] = 3'd7;
    mem[543] = 3'd0;
    mem[544] = 3'd0;
    mem[545] = 3'd7;
    mem[546] = 3'd7;
    mem[547] = 3'd7;
    mem[548] = 3'd7;
    mem[549] = 3'd7;
    mem[550] = 3'd7;
    mem[551] = 3'd7;
    mem[552] = 3'd7;
    mem[553] = 3'd0;
    mem[554] = 3'd0;
    mem[555] = 3'd0;
    mem[556] = 3'd0;
    mem[557] = 3'd7;
    mem[558] = 3'd7;
    mem[559] = 3'd0;
    mem[560] = 3'd0;
    mem[561] = 3'd7;
    mem[562] = 3'd7;
    mem[563] = 3'd7;
    mem[564] = 3'd7;
    mem[565] = 3'd7;
    mem[566] = 3'd7;
    mem[567] = 3'd7;
    mem[568] = 3'd7;
    mem[569] = 3'd0;
    mem[570] = 3'd0;
    mem[571] = 3'd0;
    mem[572] = 3'd0;
    mem[573] = 3'd7;
    mem[574] = 3'd7;
    mem[575] = 3'd0;
    mem[576] = 3'd7;
    mem[577] = 3'd7;
    mem[578] = 3'd7;
    mem[579] = 3'd7;
    mem[580] = 3'd7;
    mem[581] = 3'd7;
    mem[582] = 3'd7;
    mem[583] = 3'd7;
    mem[584] = 3'd7;
    mem[585] = 3'd0;
    mem[586] = 3'd0;
    mem[587] = 3'd0;
    mem[588] = 3'd0;
    mem[589] = 3'd7;
    mem[590] = 3'd7;
    mem[591] = 3'd0;
    mem[592] = 3'd7;
    mem[593] = 3'd7;
    mem[594] = 3'd7;
    mem[595] = 3'd7;
    mem[596] = 3'd7;
    mem[597] = 3'd7;
    mem[598] = 3'd7;
    mem[599] = 3'd7;
    mem[600] = 3'd7;
    mem[601] = 3'd0;
    mem[602] = 3'd0;
    mem[603] = 3'd0;
    mem[604] = 3'd0;
    mem[605] = 3'd7;
    mem[606] = 3'd7;
    mem[607] = 3'd0;
    mem[608] = 3'd7;
    mem[609] = 3'd7;
    mem[610] = 3'd7;
    mem[611] = 3'd7;
    mem[612] = 3'd7;
    mem[613] = 3'd7;
    mem[614] = 3'd7;
    mem[615] = 3'd7;
    mem[616] = 3'd7;
    mem[617] = 3'd0;
    mem[618] = 3'd0;
    mem[619] = 3'd0;
    mem[620] = 3'd0;
    mem[621] = 3'd7;
    mem[622] = 3'd7;
    mem[623] = 3'd0;
    mem[624] = 3'd7;
    mem[625] = 3'd7;
    mem[626] = 3'd7;
    mem[627] = 3'd7;
    mem[628] = 3'd7;
    mem[629] = 3'd7;
    mem[630] = 3'd7;
    mem[631] = 3'd7;
    mem[632] = 3'd7;
    mem[633] = 3'd0;
    mem[634] = 3'd0;
    mem[635] = 3'd0;
    mem[636] = 3'd0;
    mem[637] = 3'd7;
    mem[638] = 3'd7;
    mem[639] = 3'd0;
    mem[640] = 3'd7;
    mem[641] = 3'd7;
    mem[642] = 3'd7;
    mem[643] = 3'd7;
    mem[644] = 3'd7;
    mem[645] = 3'd7;
    mem[646] = 3'd7;
    mem[647] = 3'd7;
    mem[648] = 3'd7;
    mem[649] = 3'd0;
    mem[650] = 3'd0;
    mem[651] = 3'd0;
    mem[652] = 3'd0;
    mem[653] = 3'd7;
    mem[654] = 3'd7;
    mem[655] = 3'd0;
    mem[656] = 3'd7;
    mem[657] = 3'd7;
    mem[658] = 3'd7;
    mem[659] = 3'd7;
    mem[660] = 3'd7;
    mem[661] = 3'd7;
    mem[662] = 3'd7;
    mem[663] = 3'd7;
    mem[664] = 3'd7;
    mem[665] = 3'd0;
    mem[666] = 3'd0;
    mem[667] = 3'd0;
    mem[668] = 3'd0;
    mem[669] = 3'd7;
    mem[670] = 3'd7;
    mem[671] = 3'd0;
    mem[672] = 3'd7;
    mem[673] = 3'd7;
    mem[674] = 3'd7;
    mem[675] = 3'd7;
    mem[676] = 3'd7;
    mem[677] = 3'd7;
    mem[678] = 3'd7;
    mem[679] = 3'd7;
    mem[680] = 3'd7;
    mem[681] = 3'd0;
    mem[682] = 3'd0;
    mem[683] = 3'd0;
    mem[684] = 3'd0;
    mem[685] = 3'd0;
    mem[686] = 3'd7;
    mem[687] = 3'd0;
    mem[688] = 3'd7;
    mem[689] = 3'd7;
    mem[690] = 3'd7;
    mem[691] = 3'd7;
    mem[692] = 3'd7;
    mem[693] = 3'd7;
    mem[694] = 3'd7;
    mem[695] = 3'd7;
    mem[696] = 3'd7;
    mem[697] = 3'd0;
    mem[698] = 3'd0;
    mem[699] = 3'd0;
    mem[700] = 3'd0;
    mem[701] = 3'd0;
    mem[702] = 3'd7;
    mem[703] = 3'd0;
    mem[704] = 3'd7;
    mem[705] = 3'd7;
    mem[706] = 3'd7;
    mem[707] = 3'd7;
    mem[708] = 3'd7;
    mem[709] = 3'd7;
    mem[710] = 3'd7;
    mem[711] = 3'd7;
    mem[712] = 3'd7;
    mem[713] = 3'd0;
    mem[714] = 3'd0;
    mem[715] = 3'd0;
    mem[716] = 3'd0;
    mem[717] = 3'd0;
    mem[718] = 3'd7;
    mem[719] = 3'd0;
    mem[720] = 3'd0;
    mem[721] = 3'd0;
    mem[722] = 3'd0;
    mem[723] = 3'd0;
    mem[724] = 3'd7;
    mem[725] = 3'd7;
    mem[726] = 3'd7;
    mem[727] = 3'd0;
    mem[728] = 3'd0;
    mem[729] = 3'd0;
    mem[730] = 3'd0;
    mem[731] = 3'd0;
    mem[732] = 3'd0;
    mem[733] = 3'd0;
    mem[734] = 3'd7;
    mem[735] = 3'd0;
    mem[736] = 3'd0;
    mem[737] = 3'd0;
    mem[738] = 3'd0;
    mem[739] = 3'd0;
    mem[740] = 3'd7;
    mem[741] = 3'd7;
    mem[742] = 3'd7;
    mem[743] = 3'd0;
    mem[744] = 3'd0;
    mem[745] = 3'd0;
    mem[746] = 3'd0;
    mem[747] = 3'd0;
    mem[748] = 3'd0;
    mem[749] = 3'd0;
    mem[750] = 3'd7;
    mem[751] = 3'd0;
    mem[752] = 3'd0;
    mem[753] = 3'd0;
    mem[754] = 3'd0;
    mem[755] = 3'd0;
    mem[756] = 3'd7;
    mem[757] = 3'd7;
    mem[758] = 3'd7;
    mem[759] = 3'd0;
    mem[760] = 3'd0;
    mem[761] = 3'd0;
    mem[762] = 3'd0;
    mem[763] = 3'd0;
    mem[764] = 3'd0;
    mem[765] = 3'd0;
    mem[766] = 3'd7;
    mem[767] = 3'd0;
    mem[768] = 3'd0;
    mem[769] = 3'd0;
    mem[770] = 3'd0;
    mem[771] = 3'd0;
    mem[772] = 3'd7;
    mem[773] = 3'd7;
    mem[774] = 3'd7;
    mem[775] = 3'd0;
    mem[776] = 3'd0;
    mem[777] = 3'd0;
    mem[778] = 3'd0;
    mem[779] = 3'd0;
    mem[780] = 3'd0;
    mem[781] = 3'd0;
    mem[782] = 3'd7;
    mem[783] = 3'd0;
    mem[784] = 3'd0;
    mem[785] = 3'd0;
    mem[786] = 3'd0;
    mem[787] = 3'd0;
    mem[788] = 3'd7;
    mem[789] = 3'd7;
    mem[790] = 3'd7;
    mem[791] = 3'd0;
    mem[792] = 3'd0;
    mem[793] = 3'd0;
    mem[794] = 3'd0;
    mem[795] = 3'd0;
    mem[796] = 3'd0;
    mem[797] = 3'd0;
    mem[798] = 3'd7;
    mem[799] = 3'd0;
    mem[800] = 3'd7;
    mem[801] = 3'd0;
    mem[802] = 3'd0;
    mem[803] = 3'd0;
    mem[804] = 3'd7;
    mem[805] = 3'd7;
    mem[806] = 3'd7;
    mem[807] = 3'd0;
    mem[808] = 3'd0;
    mem[809] = 3'd0;
    mem[810] = 3'd0;
    mem[811] = 3'd0;
    mem[812] = 3'd0;
    mem[813] = 3'd0;
    mem[814] = 3'd7;
    mem[815] = 3'd0;
    mem[816] = 3'd7;
    mem[817] = 3'd0;
    mem[818] = 3'd0;
    mem[819] = 3'd0;
    mem[820] = 3'd7;
    mem[821] = 3'd7;
    mem[822] = 3'd7;
    mem[823] = 3'd0;
    mem[824] = 3'd0;
    mem[825] = 3'd0;
    mem[826] = 3'd0;
    mem[827] = 3'd0;
    mem[828] = 3'd0;
    mem[829] = 3'd0;
    mem[830] = 3'd7;
    mem[831] = 3'd0;
    mem[832] = 3'd7;
    mem[833] = 3'd0;
    mem[834] = 3'd0;
    mem[835] = 3'd0;
    mem[836] = 3'd7;
    mem[837] = 3'd7;
    mem[838] = 3'd7;
    mem[839] = 3'd0;
    mem[840] = 3'd0;
    mem[841] = 3'd0;
    mem[842] = 3'd0;
    mem[843] = 3'd0;
    mem[844] = 3'd0;
    mem[845] = 3'd0;
    mem[846] = 3'd7;
    mem[847] = 3'd0;
    mem[848] = 3'd7;
    mem[849] = 3'd0;
    mem[850] = 3'd0;
    mem[851] = 3'd0;
    mem[852] = 3'd7;
    mem[853] = 3'd7;
    mem[854] = 3'd7;
    mem[855] = 3'd0;
    mem[856] = 3'd0;
    mem[857] = 3'd0;
    mem[858] = 3'd0;
    mem[859] = 3'd0;
    mem[860] = 3'd0;
    mem[861] = 3'd0;
    mem[862] = 3'd7;
    mem[863] = 3'd0;
    mem[864] = 3'd7;
    mem[865] = 3'd0;
    mem[866] = 3'd0;
    mem[867] = 3'd0;
    mem[868] = 3'd7;
    mem[869] = 3'd7;
    mem[870] = 3'd7;
    mem[871] = 3'd0;
    mem[872] = 3'd0;
    mem[873] = 3'd0;
    mem[874] = 3'd0;
    mem[875] = 3'd0;
    mem[876] = 3'd0;
    mem[877] = 3'd0;
    mem[878] = 3'd7;
    mem[879] = 3'd0;
    mem[880] = 3'd7;
    mem[881] = 3'd0;
    mem[882] = 3'd0;
    mem[883] = 3'd0;
    mem[884] = 3'd7;
    mem[885] = 3'd7;
    mem[886] = 3'd7;
    mem[887] = 3'd0;
    mem[888] = 3'd0;
    mem[889] = 3'd0;
    mem[890] = 3'd0;
    mem[891] = 3'd0;
    mem[892] = 3'd0;
    mem[893] = 3'd0;
    mem[894] = 3'd7;
    mem[895] = 3'd7;
    mem[896] = 3'd7;
    mem[897] = 3'd0;
    mem[898] = 3'd0;
    mem[899] = 3'd0;
    mem[900] = 3'd7;
    mem[901] = 3'd7;
    mem[902] = 3'd7;
    mem[903] = 3'd0;
    mem[904] = 3'd0;
    mem[905] = 3'd0;
    mem[906] = 3'd0;
    mem[907] = 3'd0;
    mem[908] = 3'd0;
    mem[909] = 3'd0;
    mem[910] = 3'd7;
    mem[911] = 3'd7;
    mem[912] = 3'd7;
    mem[913] = 3'd0;
    mem[914] = 3'd0;
    mem[915] = 3'd0;
    mem[916] = 3'd7;
    mem[917] = 3'd7;
    mem[918] = 3'd7;
    mem[919] = 3'd0;
    mem[920] = 3'd0;
    mem[921] = 3'd0;
    mem[922] = 3'd0;
    mem[923] = 3'd0;
    mem[924] = 3'd0;
    mem[925] = 3'd0;
    mem[926] = 3'd7;
    mem[927] = 3'd7;
    mem[928] = 3'd7;
    mem[929] = 3'd0;
    mem[930] = 3'd0;
    mem[931] = 3'd0;
    mem[932] = 3'd7;
    mem[933] = 3'd7;
    mem[934] = 3'd7;
    mem[935] = 3'd7;
    mem[936] = 3'd7;
    mem[937] = 3'd7;
    mem[938] = 3'd7;
    mem[939] = 3'd7;
    mem[940] = 3'd7;
    mem[941] = 3'd0;
    mem[942] = 3'd7;
    mem[943] = 3'd7;
    mem[944] = 3'd7;
    mem[945] = 3'd0;
    mem[946] = 3'd0;
    mem[947] = 3'd0;
    mem[948] = 3'd7;
    mem[949] = 3'd7;
    mem[950] = 3'd7;
    mem[951] = 3'd7;
    mem[952] = 3'd7;
    mem[953] = 3'd7;
    mem[954] = 3'd7;
    mem[955] = 3'd7;
    mem[956] = 3'd7;
    mem[957] = 3'd0;
    mem[958] = 3'd7;
    mem[959] = 3'd7;
    mem[960] = 3'd7;
    mem[961] = 3'd0;
    mem[962] = 3'd0;
    mem[963] = 3'd0;
    mem[964] = 3'd7;
    mem[965] = 3'd7;
    mem[966] = 3'd7;
    mem[967] = 3'd7;
    mem[968] = 3'd7;
    mem[969] = 3'd7;
    mem[970] = 3'd7;
    mem[971] = 3'd7;
    mem[972] = 3'd7;
    mem[973] = 3'd0;
    mem[974] = 3'd7;
    mem[975] = 3'd7;
    mem[976] = 3'd7;
    mem[977] = 3'd0;
    mem[978] = 3'd0;
    mem[979] = 3'd0;
    mem[980] = 3'd7;
    mem[981] = 3'd7;
    mem[982] = 3'd7;
    mem[983] = 3'd7;
    mem[984] = 3'd7;
    mem[985] = 3'd7;
    mem[986] = 3'd7;
    mem[987] = 3'd7;
    mem[988] = 3'd7;
    mem[989] = 3'd0;
    mem[990] = 3'd7;
    mem[991] = 3'd7;
    mem[992] = 3'd7;
    mem[993] = 3'd0;
    mem[994] = 3'd0;
    mem[995] = 3'd0;
    mem[996] = 3'd7;
    mem[997] = 3'd7;
    mem[998] = 3'd7;
    mem[999] = 3'd7;
    mem[1000] = 3'd7;
    mem[1001] = 3'd7;
    mem[1002] = 3'd7;
    mem[1003] = 3'd7;
    mem[1004] = 3'd7;
    mem[1005] = 3'd0;
    mem[1006] = 3'd7;
    mem[1007] = 3'd7;
    mem[1008] = 3'd7;
    mem[1009] = 3'd0;
    mem[1010] = 3'd0;
    mem[1011] = 3'd0;
    mem[1012] = 3'd7;
    mem[1013] = 3'd7;
    mem[1014] = 3'd7;
    mem[1015] = 3'd7;
    mem[1016] = 3'd7;
    mem[1017] = 3'd7;
    mem[1018] = 3'd7;
    mem[1019] = 3'd7;
    mem[1020] = 3'd7;
    mem[1021] = 3'd0;
    mem[1022] = 3'd7;
    mem[1023] = 3'd7;
    mem[1024] = 3'd7;
    mem[1025] = 3'd0;
    mem[1026] = 3'd0;
    mem[1027] = 3'd0;
    mem[1028] = 3'd7;
    mem[1029] = 3'd7;
    mem[1030] = 3'd7;
    mem[1031] = 3'd7;
    mem[1032] = 3'd7;
    mem[1033] = 3'd7;
    mem[1034] = 3'd7;
    mem[1035] = 3'd7;
    mem[1036] = 3'd7;
    mem[1037] = 3'd0;
    mem[1038] = 3'd7;
    mem[1039] = 3'd7;
    mem[1040] = 3'd7;
    mem[1041] = 3'd0;
    mem[1042] = 3'd0;
    mem[1043] = 3'd0;
    mem[1044] = 3'd7;
    mem[1045] = 3'd7;
    mem[1046] = 3'd7;
    mem[1047] = 3'd7;
    mem[1048] = 3'd7;
    mem[1049] = 3'd7;
    mem[1050] = 3'd7;
    mem[1051] = 3'd7;
    mem[1052] = 3'd7;
    mem[1053] = 3'd0;
    mem[1054] = 3'd7;
    mem[1055] = 3'd7;
    mem[1056] = 3'd7;
    mem[1057] = 3'd0;
    mem[1058] = 3'd0;
    mem[1059] = 3'd0;
    mem[1060] = 3'd7;
    mem[1061] = 3'd7;
    mem[1062] = 3'd7;
    mem[1063] = 3'd7;
    mem[1064] = 3'd7;
    mem[1065] = 3'd7;
    mem[1066] = 3'd7;
    mem[1067] = 3'd7;
    mem[1068] = 3'd7;
    mem[1069] = 3'd0;
    mem[1070] = 3'd7;
    mem[1071] = 3'd7;
    mem[1072] = 3'd7;
    mem[1073] = 3'd0;
    mem[1074] = 3'd0;
    mem[1075] = 3'd0;
    mem[1076] = 3'd7;
    mem[1077] = 3'd7;
    mem[1078] = 3'd7;
    mem[1079] = 3'd7;
    mem[1080] = 3'd7;
    mem[1081] = 3'd7;
    mem[1082] = 3'd7;
    mem[1083] = 3'd7;
    mem[1084] = 3'd7;
    mem[1085] = 3'd0;
    mem[1086] = 3'd7;
    mem[1087] = 3'd7;
    mem[1088] = 3'd7;
    mem[1089] = 3'd0;
    mem[1090] = 3'd0;
    mem[1091] = 3'd0;
    mem[1092] = 3'd7;
    mem[1093] = 3'd7;
    mem[1094] = 3'd7;
    mem[1095] = 3'd7;
    mem[1096] = 3'd7;
    mem[1097] = 3'd7;
    mem[1098] = 3'd7;
    mem[1099] = 3'd7;
    mem[1100] = 3'd7;
    mem[1101] = 3'd0;
    mem[1102] = 3'd7;
    mem[1103] = 3'd7;
    mem[1104] = 3'd7;
    mem[1105] = 3'd0;
    mem[1106] = 3'd0;
    mem[1107] = 3'd0;
    mem[1108] = 3'd7;
    mem[1109] = 3'd7;
    mem[1110] = 3'd7;
    mem[1111] = 3'd7;
    mem[1112] = 3'd7;
    mem[1113] = 3'd7;
    mem[1114] = 3'd7;
    mem[1115] = 3'd7;
    mem[1116] = 3'd7;
    mem[1117] = 3'd0;
    mem[1118] = 3'd7;
    mem[1119] = 3'd7;
    mem[1120] = 3'd7;
    mem[1121] = 3'd0;
    mem[1122] = 3'd0;
    mem[1123] = 3'd0;
    mem[1124] = 3'd7;
    mem[1125] = 3'd7;
    mem[1126] = 3'd7;
    mem[1127] = 3'd7;
    mem[1128] = 3'd7;
    mem[1129] = 3'd7;
    mem[1130] = 3'd7;
    mem[1131] = 3'd7;
    mem[1132] = 3'd7;
    mem[1133] = 3'd0;
    mem[1134] = 3'd7;
    mem[1135] = 3'd7;
    mem[1136] = 3'd7;
    mem[1137] = 3'd0;
    mem[1138] = 3'd0;
    mem[1139] = 3'd0;
    mem[1140] = 3'd7;
    mem[1141] = 3'd7;
    mem[1142] = 3'd7;
    mem[1143] = 3'd7;
    mem[1144] = 3'd7;
    mem[1145] = 3'd7;
    mem[1146] = 3'd7;
    mem[1147] = 3'd7;
    mem[1148] = 3'd7;
    mem[1149] = 3'd0;
    mem[1150] = 3'd7;
    mem[1151] = 3'd7;
    mem[1152] = 3'd7;
    mem[1153] = 3'd0;
    mem[1154] = 3'd0;
    mem[1155] = 3'd0;
    mem[1156] = 3'd7;
    mem[1157] = 3'd7;
    mem[1158] = 3'd7;
    mem[1159] = 3'd7;
    mem[1160] = 3'd7;
    mem[1161] = 3'd7;
    mem[1162] = 3'd7;
    mem[1163] = 3'd7;
    mem[1164] = 3'd7;
    mem[1165] = 3'd0;
    mem[1166] = 3'd7;
    mem[1167] = 3'd7;
    mem[1168] = 3'd7;
    mem[1169] = 3'd0;
    mem[1170] = 3'd0;
    mem[1171] = 3'd0;
    mem[1172] = 3'd7;
    mem[1173] = 3'd7;
    mem[1174] = 3'd7;
    mem[1175] = 3'd7;
    mem[1176] = 3'd7;
    mem[1177] = 3'd7;
    mem[1178] = 3'd7;
    mem[1179] = 3'd7;
    mem[1180] = 3'd7;
    mem[1181] = 3'd0;
    mem[1182] = 3'd7;
    mem[1183] = 3'd0;
    mem[1184] = 3'd7;
    mem[1185] = 3'd0;
    mem[1186] = 3'd0;
    mem[1187] = 3'd0;
    mem[1188] = 3'd7;
    mem[1189] = 3'd7;
    mem[1190] = 3'd7;
    mem[1191] = 3'd7;
    mem[1192] = 3'd7;
    mem[1193] = 3'd7;
    mem[1194] = 3'd7;
    mem[1195] = 3'd7;
    mem[1196] = 3'd7;
    mem[1197] = 3'd0;
    mem[1198] = 3'd7;
    mem[1199] = 3'd0;
    mem[1200] = 3'd7;
    mem[1201] = 3'd0;
    mem[1202] = 3'd0;
    mem[1203] = 3'd0;
    mem[1204] = 3'd7;
    mem[1205] = 3'd7;
    mem[1206] = 3'd7;
    mem[1207] = 3'd7;
    mem[1208] = 3'd7;
    mem[1209] = 3'd7;
    mem[1210] = 3'd7;
    mem[1211] = 3'd7;
    mem[1212] = 3'd7;
    mem[1213] = 3'd0;
    mem[1214] = 3'd7;
    mem[1215] = 3'd0;
    mem[1216] = 3'd7;
    mem[1217] = 3'd0;
    mem[1218] = 3'd0;
    mem[1219] = 3'd0;
    mem[1220] = 3'd7;
    mem[1221] = 3'd7;
    mem[1222] = 3'd7;
    mem[1223] = 3'd0;
    mem[1224] = 3'd7;
    mem[1225] = 3'd7;
    mem[1226] = 3'd7;
    mem[1227] = 3'd0;
    mem[1228] = 3'd0;
    mem[1229] = 3'd0;
    mem[1230] = 3'd7;
    mem[1231] = 3'd0;
    mem[1232] = 3'd7;
    mem[1233] = 3'd0;
    mem[1234] = 3'd0;
    mem[1235] = 3'd0;
    mem[1236] = 3'd7;
    mem[1237] = 3'd7;
    mem[1238] = 3'd7;
    mem[1239] = 3'd0;
    mem[1240] = 3'd7;
    mem[1241] = 3'd7;
    mem[1242] = 3'd7;
    mem[1243] = 3'd0;
    mem[1244] = 3'd0;
    mem[1245] = 3'd0;
    mem[1246] = 3'd7;
    mem[1247] = 3'd0;
    mem[1248] = 3'd7;
    mem[1249] = 3'd0;
    mem[1250] = 3'd0;
    mem[1251] = 3'd0;
    mem[1252] = 3'd7;
    mem[1253] = 3'd7;
    mem[1254] = 3'd7;
    mem[1255] = 3'd0;
    mem[1256] = 3'd7;
    mem[1257] = 3'd7;
    mem[1258] = 3'd7;
    mem[1259] = 3'd0;
    mem[1260] = 3'd0;
    mem[1261] = 3'd0;
    mem[1262] = 3'd7;
    mem[1263] = 3'd0;
    mem[1264] = 3'd7;
    mem[1265] = 3'd0;
    mem[1266] = 3'd0;
    mem[1267] = 3'd0;
    mem[1268] = 3'd7;
    mem[1269] = 3'd7;
    mem[1270] = 3'd7;
    mem[1271] = 3'd0;
    mem[1272] = 3'd7;
    mem[1273] = 3'd7;
    mem[1274] = 3'd7;
    mem[1275] = 3'd0;
    mem[1276] = 3'd0;
    mem[1277] = 3'd0;
    mem[1278] = 3'd7;
    mem[1279] = 3'd0;
    mem[1280] = 3'd7;
    mem[1281] = 3'd0;
    mem[1282] = 3'd0;
    mem[1283] = 3'd0;
    mem[1284] = 3'd7;
    mem[1285] = 3'd7;
    mem[1286] = 3'd7;
    mem[1287] = 3'd0;
    mem[1288] = 3'd7;
    mem[1289] = 3'd7;
    mem[1290] = 3'd7;
    mem[1291] = 3'd0;
    mem[1292] = 3'd0;
    mem[1293] = 3'd0;
    mem[1294] = 3'd7;
    mem[1295] = 3'd0;
    mem[1296] = 3'd7;
    mem[1297] = 3'd7;
    mem[1298] = 3'd0;
    mem[1299] = 3'd0;
    mem[1300] = 3'd7;
    mem[1301] = 3'd7;
    mem[1302] = 3'd7;
    mem[1303] = 3'd0;
    mem[1304] = 3'd7;
    mem[1305] = 3'd7;
    mem[1306] = 3'd7;
    mem[1307] = 3'd0;
    mem[1308] = 3'd0;
    mem[1309] = 3'd0;
    mem[1310] = 3'd7;
    mem[1311] = 3'd0;
    mem[1312] = 3'd7;
    mem[1313] = 3'd7;
    mem[1314] = 3'd0;
    mem[1315] = 3'd0;
    mem[1316] = 3'd7;
    mem[1317] = 3'd7;
    mem[1318] = 3'd7;
    mem[1319] = 3'd0;
    mem[1320] = 3'd7;
    mem[1321] = 3'd7;
    mem[1322] = 3'd7;
    mem[1323] = 3'd0;
    mem[1324] = 3'd0;
    mem[1325] = 3'd0;
    mem[1326] = 3'd7;
    mem[1327] = 3'd0;
    mem[1328] = 3'd7;
    mem[1329] = 3'd7;
    mem[1330] = 3'd0;
    mem[1331] = 3'd0;
    mem[1332] = 3'd7;
    mem[1333] = 3'd7;
    mem[1334] = 3'd7;
    mem[1335] = 3'd0;
    mem[1336] = 3'd7;
    mem[1337] = 3'd7;
    mem[1338] = 3'd7;
    mem[1339] = 3'd0;
    mem[1340] = 3'd0;
    mem[1341] = 3'd0;
    mem[1342] = 3'd7;
    mem[1343] = 3'd0;
    mem[1344] = 3'd7;
    mem[1345] = 3'd7;
    mem[1346] = 3'd0;
    mem[1347] = 3'd0;
    mem[1348] = 3'd7;
    mem[1349] = 3'd7;
    mem[1350] = 3'd7;
    mem[1351] = 3'd0;
    mem[1352] = 3'd7;
    mem[1353] = 3'd7;
    mem[1354] = 3'd7;
    mem[1355] = 3'd0;
    mem[1356] = 3'd0;
    mem[1357] = 3'd0;
    mem[1358] = 3'd7;
    mem[1359] = 3'd0;
    mem[1360] = 3'd7;
    mem[1361] = 3'd7;
    mem[1362] = 3'd0;
    mem[1363] = 3'd0;
    mem[1364] = 3'd7;
    mem[1365] = 3'd7;
    mem[1366] = 3'd7;
    mem[1367] = 3'd0;
    mem[1368] = 3'd7;
    mem[1369] = 3'd7;
    mem[1370] = 3'd7;
    mem[1371] = 3'd0;
    mem[1372] = 3'd0;
    mem[1373] = 3'd0;
    mem[1374] = 3'd7;
    mem[1375] = 3'd0;
    mem[1376] = 3'd7;
    mem[1377] = 3'd7;
    mem[1378] = 3'd0;
    mem[1379] = 3'd0;
    mem[1380] = 3'd7;
    mem[1381] = 3'd7;
    mem[1382] = 3'd7;
    mem[1383] = 3'd0;
    mem[1384] = 3'd7;
    mem[1385] = 3'd7;
    mem[1386] = 3'd7;
    mem[1387] = 3'd0;
    mem[1388] = 3'd0;
    mem[1389] = 3'd7;
    mem[1390] = 3'd7;
    mem[1391] = 3'd0;
    mem[1392] = 3'd7;
    mem[1393] = 3'd7;
    mem[1394] = 3'd0;
    mem[1395] = 3'd0;
    mem[1396] = 3'd0;
    mem[1397] = 3'd0;
    mem[1398] = 3'd0;
    mem[1399] = 3'd0;
    mem[1400] = 3'd7;
    mem[1401] = 3'd7;
    mem[1402] = 3'd7;
    mem[1403] = 3'd0;
    mem[1404] = 3'd0;
    mem[1405] = 3'd7;
    mem[1406] = 3'd7;
    mem[1407] = 3'd0;
    mem[1408] = 3'd7;
    mem[1409] = 3'd7;
    mem[1410] = 3'd0;
    mem[1411] = 3'd0;
    mem[1412] = 3'd0;
    mem[1413] = 3'd0;
    mem[1414] = 3'd0;
    mem[1415] = 3'd0;
    mem[1416] = 3'd7;
    mem[1417] = 3'd7;
    mem[1418] = 3'd7;
    mem[1419] = 3'd0;
    mem[1420] = 3'd0;
    mem[1421] = 3'd7;
    mem[1422] = 3'd7;
    mem[1423] = 3'd0;
    mem[1424] = 3'd7;
    mem[1425] = 3'd7;
    mem[1426] = 3'd0;
    mem[1427] = 3'd0;
    mem[1428] = 3'd0;
    mem[1429] = 3'd0;
    mem[1430] = 3'd0;
    mem[1431] = 3'd0;
    mem[1432] = 3'd7;
    mem[1433] = 3'd7;
    mem[1434] = 3'd7;
    mem[1435] = 3'd0;
    mem[1436] = 3'd0;
    mem[1437] = 3'd7;
    mem[1438] = 3'd7;
    mem[1439] = 3'd0;
    mem[1440] = 3'd7;
    mem[1441] = 3'd7;
    mem[1442] = 3'd0;
    mem[1443] = 3'd0;
    mem[1444] = 3'd0;
    mem[1445] = 3'd0;
    mem[1446] = 3'd0;
    mem[1447] = 3'd0;
    mem[1448] = 3'd7;
    mem[1449] = 3'd7;
    mem[1450] = 3'd7;
    mem[1451] = 3'd0;
    mem[1452] = 3'd0;
    mem[1453] = 3'd7;
    mem[1454] = 3'd7;
    mem[1455] = 3'd0;
    mem[1456] = 3'd7;
    mem[1457] = 3'd7;
    mem[1458] = 3'd0;
    mem[1459] = 3'd0;
    mem[1460] = 3'd0;
    mem[1461] = 3'd0;
    mem[1462] = 3'd0;
    mem[1463] = 3'd0;
    mem[1464] = 3'd7;
    mem[1465] = 3'd7;
    mem[1466] = 3'd7;
    mem[1467] = 3'd0;
    mem[1468] = 3'd0;
    mem[1469] = 3'd7;
    mem[1470] = 3'd7;
    mem[1471] = 3'd0;
    mem[1472] = 3'd0;
    mem[1473] = 3'd7;
    mem[1474] = 3'd0;
    mem[1475] = 3'd0;
    mem[1476] = 3'd0;
    mem[1477] = 3'd0;
    mem[1478] = 3'd0;
    mem[1479] = 3'd0;
    mem[1480] = 3'd7;
    mem[1481] = 3'd7;
    mem[1482] = 3'd7;
    mem[1483] = 3'd0;
    mem[1484] = 3'd0;
    mem[1485] = 3'd7;
    mem[1486] = 3'd7;
    mem[1487] = 3'd0;
    mem[1488] = 3'd0;
    mem[1489] = 3'd7;
    mem[1490] = 3'd0;
    mem[1491] = 3'd0;
    mem[1492] = 3'd0;
    mem[1493] = 3'd0;
    mem[1494] = 3'd0;
    mem[1495] = 3'd0;
    mem[1496] = 3'd7;
    mem[1497] = 3'd7;
    mem[1498] = 3'd7;
    mem[1499] = 3'd0;
    mem[1500] = 3'd0;
    mem[1501] = 3'd7;
    mem[1502] = 3'd7;
    mem[1503] = 3'd0;
    mem[1504] = 3'd0;
    mem[1505] = 3'd7;
    mem[1506] = 3'd0;
    mem[1507] = 3'd0;
    mem[1508] = 3'd0;
    mem[1509] = 3'd0;
    mem[1510] = 3'd0;
    mem[1511] = 3'd0;
    mem[1512] = 3'd7;
    mem[1513] = 3'd7;
    mem[1514] = 3'd7;
    mem[1515] = 3'd0;
    mem[1516] = 3'd0;
    mem[1517] = 3'd7;
    mem[1518] = 3'd7;
    mem[1519] = 3'd0;
    mem[1520] = 3'd0;
    mem[1521] = 3'd7;
    mem[1522] = 3'd0;
    mem[1523] = 3'd0;
    mem[1524] = 3'd0;
    mem[1525] = 3'd0;
    mem[1526] = 3'd0;
    mem[1527] = 3'd0;
    mem[1528] = 3'd7;
    mem[1529] = 3'd7;
    mem[1530] = 3'd7;
    mem[1531] = 3'd0;
    mem[1532] = 3'd0;
    mem[1533] = 3'd7;
    mem[1534] = 3'd7;
    mem[1535] = 3'd0;
    mem[1536] = 3'd0;
    mem[1537] = 3'd7;
    mem[1538] = 3'd7;
    mem[1539] = 3'd0;
    mem[1540] = 3'd0;
    mem[1541] = 3'd0;
    mem[1542] = 3'd0;
    mem[1543] = 3'd0;
    mem[1544] = 3'd7;
    mem[1545] = 3'd7;
    mem[1546] = 3'd7;
    mem[1547] = 3'd0;
    mem[1548] = 3'd0;
    mem[1549] = 3'd7;
    mem[1550] = 3'd0;
    mem[1551] = 3'd0;
    mem[1552] = 3'd0;
    mem[1553] = 3'd7;
    mem[1554] = 3'd7;
    mem[1555] = 3'd0;
    mem[1556] = 3'd0;
    mem[1557] = 3'd0;
    mem[1558] = 3'd0;
    mem[1559] = 3'd0;
    mem[1560] = 3'd7;
    mem[1561] = 3'd7;
    mem[1562] = 3'd7;
    mem[1563] = 3'd0;
    mem[1564] = 3'd0;
    mem[1565] = 3'd7;
    mem[1566] = 3'd0;
    mem[1567] = 3'd0;
    mem[1568] = 3'd0;
    mem[1569] = 3'd7;
    mem[1570] = 3'd7;
    mem[1571] = 3'd0;
    mem[1572] = 3'd0;
    mem[1573] = 3'd0;
    mem[1574] = 3'd0;
    mem[1575] = 3'd0;
    mem[1576] = 3'd7;
    mem[1577] = 3'd7;
    mem[1578] = 3'd7;
    mem[1579] = 3'd0;
    mem[1580] = 3'd7;
    mem[1581] = 3'd7;
    mem[1582] = 3'd0;
    mem[1583] = 3'd0;
    mem[1584] = 3'd0;
    mem[1585] = 3'd7;
    mem[1586] = 3'd7;
    mem[1587] = 3'd0;
    mem[1588] = 3'd0;
    mem[1589] = 3'd0;
    mem[1590] = 3'd0;
    mem[1591] = 3'd0;
    mem[1592] = 3'd7;
    mem[1593] = 3'd7;
    mem[1594] = 3'd7;
    mem[1595] = 3'd0;
    mem[1596] = 3'd7;
    mem[1597] = 3'd7;
    mem[1598] = 3'd0;
    mem[1599] = 3'd0;
    mem[1600] = 3'd0;
    mem[1601] = 3'd7;
    mem[1602] = 3'd7;
    mem[1603] = 3'd0;
    mem[1604] = 3'd0;
    mem[1605] = 3'd0;
    mem[1606] = 3'd0;
    mem[1607] = 3'd0;
    mem[1608] = 3'd7;
    mem[1609] = 3'd7;
    mem[1610] = 3'd7;
    mem[1611] = 3'd0;
    mem[1612] = 3'd7;
    mem[1613] = 3'd7;
    mem[1614] = 3'd0;
    mem[1615] = 3'd0;
    mem[1616] = 3'd0;
    mem[1617] = 3'd7;
    mem[1618] = 3'd7;
    mem[1619] = 3'd0;
    mem[1620] = 3'd0;
    mem[1621] = 3'd0;
    mem[1622] = 3'd0;
    mem[1623] = 3'd0;
    mem[1624] = 3'd7;
    mem[1625] = 3'd7;
    mem[1626] = 3'd7;
    mem[1627] = 3'd0;
    mem[1628] = 3'd7;
    mem[1629] = 3'd7;
    mem[1630] = 3'd0;
    mem[1631] = 3'd0;
    mem[1632] = 3'd0;
    mem[1633] = 3'd7;
    mem[1634] = 3'd7;
    mem[1635] = 3'd0;
    mem[1636] = 3'd0;
    mem[1637] = 3'd0;
    mem[1638] = 3'd0;
    mem[1639] = 3'd0;
    mem[1640] = 3'd7;
    mem[1641] = 3'd7;
    mem[1642] = 3'd7;
    mem[1643] = 3'd0;
    mem[1644] = 3'd7;
    mem[1645] = 3'd7;
    mem[1646] = 3'd0;
    mem[1647] = 3'd0;
    mem[1648] = 3'd0;
    mem[1649] = 3'd7;
    mem[1650] = 3'd7;
    mem[1651] = 3'd0;
    mem[1652] = 3'd0;
    mem[1653] = 3'd0;
    mem[1654] = 3'd0;
    mem[1655] = 3'd0;
    mem[1656] = 3'd7;
    mem[1657] = 3'd7;
    mem[1658] = 3'd7;
    mem[1659] = 3'd0;
    mem[1660] = 3'd7;
    mem[1661] = 3'd7;
    mem[1662] = 3'd0;
    mem[1663] = 3'd0;
    mem[1664] = 3'd0;
    mem[1665] = 3'd7;
    mem[1666] = 3'd7;
    mem[1667] = 3'd7;
    mem[1668] = 3'd0;
    mem[1669] = 3'd0;
    mem[1670] = 3'd0;
    mem[1671] = 3'd0;
    mem[1672] = 3'd7;
    mem[1673] = 3'd7;
    mem[1674] = 3'd7;
    mem[1675] = 3'd0;
    mem[1676] = 3'd7;
    mem[1677] = 3'd7;
    mem[1678] = 3'd0;
    mem[1679] = 3'd0;
    mem[1680] = 3'd0;
    mem[1681] = 3'd0;
    mem[1682] = 3'd7;
    mem[1683] = 3'd7;
    mem[1684] = 3'd0;
    mem[1685] = 3'd0;
    mem[1686] = 3'd0;
    mem[1687] = 3'd0;
    mem[1688] = 3'd7;
    mem[1689] = 3'd7;
    mem[1690] = 3'd7;
    mem[1691] = 3'd0;
    mem[1692] = 3'd7;
    mem[1693] = 3'd7;
    mem[1694] = 3'd0;
    mem[1695] = 3'd0;
    mem[1696] = 3'd0;
    mem[1697] = 3'd0;
    mem[1698] = 3'd7;
    mem[1699] = 3'd7;
    mem[1700] = 3'd0;
    mem[1701] = 3'd0;
    mem[1702] = 3'd0;
    mem[1703] = 3'd0;
    mem[1704] = 3'd7;
    mem[1705] = 3'd7;
    mem[1706] = 3'd7;
    mem[1707] = 3'd7;
    mem[1708] = 3'd7;
    mem[1709] = 3'd7;
    mem[1710] = 3'd0;
    mem[1711] = 3'd0;
    mem[1712] = 3'd0;
    mem[1713] = 3'd0;
    mem[1714] = 3'd7;
    mem[1715] = 3'd7;
    mem[1716] = 3'd0;
    mem[1717] = 3'd0;
    mem[1718] = 3'd0;
    mem[1719] = 3'd0;
    mem[1720] = 3'd7;
    mem[1721] = 3'd7;
    mem[1722] = 3'd7;
    mem[1723] = 3'd7;
    mem[1724] = 3'd7;
    mem[1725] = 3'd0;
    mem[1726] = 3'd0;
    mem[1727] = 3'd0;
    mem[1728] = 3'd0;
    mem[1729] = 3'd0;
    mem[1730] = 3'd7;
    mem[1731] = 3'd7;
    mem[1732] = 3'd0;
    mem[1733] = 3'd0;
    mem[1734] = 3'd0;
    mem[1735] = 3'd0;
    mem[1736] = 3'd7;
    mem[1737] = 3'd7;
    mem[1738] = 3'd7;
    mem[1739] = 3'd7;
    mem[1740] = 3'd7;
    mem[1741] = 3'd0;
    mem[1742] = 3'd0;
    mem[1743] = 3'd0;
    mem[1744] = 3'd0;
    mem[1745] = 3'd0;
    mem[1746] = 3'd7;
    mem[1747] = 3'd7;
    mem[1748] = 3'd0;
    mem[1749] = 3'd0;
    mem[1750] = 3'd0;
    mem[1751] = 3'd0;
    mem[1752] = 3'd7;
    mem[1753] = 3'd7;
    mem[1754] = 3'd7;
    mem[1755] = 3'd7;
    mem[1756] = 3'd7;
    mem[1757] = 3'd0;
    mem[1758] = 3'd0;
    mem[1759] = 3'd0;
    mem[1760] = 3'd0;
    mem[1761] = 3'd0;
    mem[1762] = 3'd7;
    mem[1763] = 3'd7;
    mem[1764] = 3'd7;
    mem[1765] = 3'd0;
    mem[1766] = 3'd0;
    mem[1767] = 3'd0;
    mem[1768] = 3'd7;
    mem[1769] = 3'd7;
    mem[1770] = 3'd7;
    mem[1771] = 3'd7;
    mem[1772] = 3'd7;
    mem[1773] = 3'd0;
    mem[1774] = 3'd0;
    mem[1775] = 3'd0;
    mem[1776] = 3'd0;
    mem[1777] = 3'd0;
    mem[1778] = 3'd7;
    mem[1779] = 3'd7;
    mem[1780] = 3'd7;
    mem[1781] = 3'd0;
    mem[1782] = 3'd0;
    mem[1783] = 3'd0;
    mem[1784] = 3'd7;
    mem[1785] = 3'd7;
    mem[1786] = 3'd7;
    mem[1787] = 3'd7;
    mem[1788] = 3'd7;
    mem[1789] = 3'd0;
    mem[1790] = 3'd0;
    mem[1791] = 3'd0;
    mem[1792] = 3'd0;
    mem[1793] = 3'd0;
    mem[1794] = 3'd7;
    mem[1795] = 3'd7;
    mem[1796] = 3'd7;
    mem[1797] = 3'd0;
    mem[1798] = 3'd0;
    mem[1799] = 3'd0;
    mem[1800] = 3'd7;
    mem[1801] = 3'd7;
    mem[1802] = 3'd7;
    mem[1803] = 3'd7;
    mem[1804] = 3'd7;
    mem[1805] = 3'd0;
    mem[1806] = 3'd0;
    mem[1807] = 3'd0;
    mem[1808] = 3'd0;
    mem[1809] = 3'd0;
    mem[1810] = 3'd0;
    mem[1811] = 3'd7;
    mem[1812] = 3'd7;
    mem[1813] = 3'd7;
    mem[1814] = 3'd0;
    mem[1815] = 3'd0;
    mem[1816] = 3'd7;
    mem[1817] = 3'd7;
    mem[1818] = 3'd7;
    mem[1819] = 3'd7;
    mem[1820] = 3'd7;
    mem[1821] = 3'd0;
    mem[1822] = 3'd0;
    mem[1823] = 3'd0;
    mem[1824] = 3'd0;
    mem[1825] = 3'd0;
    mem[1826] = 3'd0;
    mem[1827] = 3'd7;
    mem[1828] = 3'd7;
    mem[1829] = 3'd7;
    mem[1830] = 3'd0;
    mem[1831] = 3'd0;
    mem[1832] = 3'd7;
    mem[1833] = 3'd7;
    mem[1834] = 3'd7;
    mem[1835] = 3'd7;
    mem[1836] = 3'd0;
    mem[1837] = 3'd0;
    mem[1838] = 3'd0;
    mem[1839] = 3'd0;
    mem[1840] = 3'd0;
    mem[1841] = 3'd0;
    mem[1842] = 3'd0;
    mem[1843] = 3'd7;
    mem[1844] = 3'd7;
    mem[1845] = 3'd7;
    mem[1846] = 3'd0;
    mem[1847] = 3'd0;
    mem[1848] = 3'd7;
    mem[1849] = 3'd7;
    mem[1850] = 3'd7;
    mem[1851] = 3'd7;
    mem[1852] = 3'd0;
    mem[1853] = 3'd0;
    mem[1854] = 3'd0;
    mem[1855] = 3'd0;
    mem[1856] = 3'd0;
    mem[1857] = 3'd0;
    mem[1858] = 3'd0;
    mem[1859] = 3'd7;
    mem[1860] = 3'd7;
    mem[1861] = 3'd7;
    mem[1862] = 3'd7;
    mem[1863] = 3'd7;
    mem[1864] = 3'd7;
    mem[1865] = 3'd7;
    mem[1866] = 3'd7;
    mem[1867] = 3'd7;
    mem[1868] = 3'd0;
    mem[1869] = 3'd0;
    mem[1870] = 3'd0;
    mem[1871] = 3'd0;
    mem[1872] = 3'd0;
    mem[1873] = 3'd0;
    mem[1874] = 3'd0;
    mem[1875] = 3'd7;
    mem[1876] = 3'd7;
    mem[1877] = 3'd7;
    mem[1878] = 3'd7;
    mem[1879] = 3'd7;
    mem[1880] = 3'd7;
    mem[1881] = 3'd7;
    mem[1882] = 3'd7;
    mem[1883] = 3'd7;
    mem[1884] = 3'd0;
    mem[1885] = 3'd0;
    mem[1886] = 3'd0;
    mem[1887] = 3'd0;
    mem[1888] = 3'd0;
    mem[1889] = 3'd0;
    mem[1890] = 3'd0;
    mem[1891] = 3'd0;
    mem[1892] = 3'd7;
    mem[1893] = 3'd7;
    mem[1894] = 3'd7;
    mem[1895] = 3'd7;
    mem[1896] = 3'd7;
    mem[1897] = 3'd7;
    mem[1898] = 3'd7;
    mem[1899] = 3'd7;
    mem[1900] = 3'd0;
    mem[1901] = 3'd0;
    mem[1902] = 3'd0;
    mem[1903] = 3'd0;
    mem[1904] = 3'd0;
    mem[1905] = 3'd0;
    mem[1906] = 3'd0;
    mem[1907] = 3'd0;
    mem[1908] = 3'd7;
    mem[1909] = 3'd7;
    mem[1910] = 3'd7;
    mem[1911] = 3'd7;
    mem[1912] = 3'd7;
    mem[1913] = 3'd7;
    mem[1914] = 3'd7;
    mem[1915] = 3'd0;
    mem[1916] = 3'd0;
    mem[1917] = 3'd0;
    mem[1918] = 3'd0;
    mem[1919] = 3'd0;
    mem[1920] = 3'd0;
    mem[1921] = 3'd0;
    mem[1922] = 3'd0;
    mem[1923] = 3'd0;
    mem[1924] = 3'd7;
    mem[1925] = 3'd7;
    mem[1926] = 3'd7;
    mem[1927] = 3'd7;
    mem[1928] = 3'd7;
    mem[1929] = 3'd7;
    mem[1930] = 3'd7;
    mem[1931] = 3'd0;
    mem[1932] = 3'd0;
    mem[1933] = 3'd0;
    mem[1934] = 3'd0;
    mem[1935] = 3'd0;
    mem[1936] = 3'd0;
    mem[1937] = 3'd0;
    mem[1938] = 3'd0;
    mem[1939] = 3'd0;
    mem[1940] = 3'd7;
    mem[1941] = 3'd7;
    mem[1942] = 3'd7;
    mem[1943] = 3'd7;
    mem[1944] = 3'd7;
    mem[1945] = 3'd7;
    mem[1946] = 3'd7;
    mem[1947] = 3'd0;
    mem[1948] = 3'd0;
    mem[1949] = 3'd0;
    mem[1950] = 3'd0;
    mem[1951] = 3'd0;
    mem[1952] = 3'd0;
    mem[1953] = 3'd0;
    mem[1954] = 3'd0;
    mem[1955] = 3'd0;
    mem[1956] = 3'd0;
    mem[1957] = 3'd7;
    mem[1958] = 3'd7;
    mem[1959] = 3'd7;
    mem[1960] = 3'd7;
    mem[1961] = 3'd7;
    mem[1962] = 3'd7;
    mem[1963] = 3'd0;
    mem[1964] = 3'd0;
    mem[1965] = 3'd0;
    mem[1966] = 3'd0;
    mem[1967] = 3'd0;
    mem[1968] = 3'd0;
    mem[1969] = 3'd0;
    mem[1970] = 3'd0;
    mem[1971] = 3'd0;
    mem[1972] = 3'd0;
    mem[1973] = 3'd7;
    mem[1974] = 3'd7;
    mem[1975] = 3'd7;
    mem[1976] = 3'd7;
    mem[1977] = 3'd7;
    mem[1978] = 3'd0;
    mem[1979] = 3'd0;
    mem[1980] = 3'd0;
    mem[1981] = 3'd0;
    mem[1982] = 3'd0;
    mem[1983] = 3'd0;
    mem[1984] = 3'd0;
    mem[1985] = 3'd0;
    mem[1986] = 3'd0;
    mem[1987] = 3'd0;
    mem[1988] = 3'd0;
    mem[1989] = 3'd7;
    mem[1990] = 3'd7;
    mem[1991] = 3'd7;
    mem[1992] = 3'd7;
    mem[1993] = 3'd7;
    mem[1994] = 3'd0;
    mem[1995] = 3'd0;
    mem[1996] = 3'd0;
    mem[1997] = 3'd0;
    mem[1998] = 3'd0;
    mem[1999] = 3'd0;
    mem[2000] = 3'd0;
    mem[2001] = 3'd0;
    mem[2002] = 3'd0;
    mem[2003] = 3'd0;
    mem[2004] = 3'd0;
    mem[2005] = 3'd0;
    mem[2006] = 3'd7;
    mem[2007] = 3'd7;
    mem[2008] = 3'd7;
    mem[2009] = 3'd0;
    mem[2010] = 3'd0;
    mem[2011] = 3'd0;
    mem[2012] = 3'd0;
    mem[2013] = 3'd0;
    mem[2014] = 3'd0;
    mem[2015] = 3'd0;
    mem[2016] = 3'd0;
    mem[2017] = 3'd0;
    mem[2018] = 3'd0;
    mem[2019] = 3'd0;
    mem[2020] = 3'd0;
    mem[2021] = 3'd0;
    mem[2022] = 3'd7;
    mem[2023] = 3'd7;
    mem[2024] = 3'd7;
    mem[2025] = 3'd0;
    mem[2026] = 3'd0;
    mem[2027] = 3'd0;
    mem[2028] = 3'd0;
    mem[2029] = 3'd0;
    mem[2030] = 3'd0;
    mem[2031] = 3'd0;
    mem[2032] = 3'd0;
    mem[2033] = 3'd0;
    mem[2034] = 3'd0;
    mem[2035] = 3'd0;
    mem[2036] = 3'd0;
    mem[2037] = 3'd0;
    mem[2038] = 3'd0;
    mem[2039] = 3'd0;
    mem[2040] = 3'd0;
    mem[2041] = 3'd0;
    mem[2042] = 3'd0;
    mem[2043] = 3'd0;
    mem[2044] = 3'd0;
    mem[2045] = 3'd0;
    mem[2046] = 3'd0;
    mem[2047] = 3'd0;
  end

    wire [10:0] addr = {y[6:0], x[6:3]};
  assign pixel[2:0] = mem[addr];

endmodule

module bitmap_rom (
    input wire [6:0] x,
    input wire [6:0] y,
    output wire red_pixel,
    output wire green_pixel,
    output wire blue_pixel
);

  reg [7:0] red_mem[2047:0];
  reg [7:0] green_mem[2047:0];
  reg [7:0] blue_mem[2047:0];
  initial begin
    red_mem[0] = 8'h00;
    red_mem[1] = 8'h00;
    red_mem[2] = 8'h00;
    red_mem[3] = 8'h00;
    red_mem[4] = 8'h00;
    red_mem[5] = 8'h00;
    red_mem[6] = 8'h00;
    red_mem[7] = 8'h00;
    red_mem[8] = 8'h00;
    red_mem[9] = 8'h00;
    red_mem[10] = 8'h00;
    red_mem[11] = 8'h00;
    red_mem[12] = 8'h00;
    red_mem[13] = 8'h00;
    red_mem[14] = 8'h00;
    red_mem[15] = 8'h00;
    red_mem[16] = 8'h00;
    red_mem[17] = 8'h00;
    red_mem[18] = 8'h00;
    red_mem[19] = 8'h00;
    red_mem[20] = 8'h00;
    red_mem[21] = 8'h00;
    red_mem[22] = 8'h00;
    red_mem[23] = 8'h00;
    red_mem[24] = 8'h00;
    red_mem[25] = 8'h00;
    red_mem[26] = 8'h00;
    red_mem[27] = 8'h00;
    red_mem[28] = 8'h00;
    red_mem[29] = 8'h00;
    red_mem[30] = 8'h00;
    red_mem[31] = 8'h00;
    red_mem[32] = 8'h00;
    red_mem[33] = 8'h00;
    red_mem[34] = 8'h00;
    red_mem[35] = 8'h00;
    red_mem[36] = 8'h00;
    red_mem[37] = 8'h00;
    red_mem[38] = 8'h00;
    red_mem[39] = 8'h00;
    red_mem[40] = 8'h00;
    red_mem[41] = 8'h00;
    red_mem[42] = 8'h00;
    red_mem[43] = 8'h00;
    red_mem[44] = 8'h00;
    red_mem[45] = 8'h00;
    red_mem[46] = 8'h00;
    red_mem[47] = 8'h00;
    red_mem[48] = 8'h00;
    red_mem[49] = 8'h00;
    red_mem[50] = 8'h00;
    red_mem[51] = 8'h00;
    red_mem[52] = 8'h00;
    red_mem[53] = 8'h00;
    red_mem[54] = 8'h00;
    red_mem[55] = 8'h00;
    red_mem[56] = 8'h00;
    red_mem[57] = 8'h00;
    red_mem[58] = 8'h00;
    red_mem[59] = 8'h00;
    red_mem[60] = 8'h00;
    red_mem[61] = 8'h00;
    red_mem[62] = 8'h00;
    red_mem[63] = 8'h00;
    red_mem[64] = 8'h00;
    red_mem[65] = 8'h00;
    red_mem[66] = 8'h00;
    red_mem[67] = 8'h00;
    red_mem[68] = 8'h00;
    red_mem[69] = 8'h00;
    red_mem[70] = 8'h00;
    red_mem[71] = 8'h00;
    red_mem[72] = 8'h00;
    red_mem[73] = 8'h00;
    red_mem[74] = 8'h00;
    red_mem[75] = 8'h00;
    red_mem[76] = 8'h00;
    red_mem[77] = 8'h00;
    red_mem[78] = 8'h00;
    red_mem[79] = 8'h00;
    red_mem[80] = 8'h00;
    red_mem[81] = 8'h00;
    red_mem[82] = 8'h00;
    red_mem[83] = 8'h00;
    red_mem[84] = 8'h00;
    red_mem[85] = 8'h00;
    red_mem[86] = 8'h00;
    red_mem[87] = 8'h00;
    red_mem[88] = 8'h00;
    red_mem[89] = 8'h00;
    red_mem[90] = 8'h00;
    red_mem[91] = 8'h00;
    red_mem[92] = 8'h00;
    red_mem[93] = 8'h00;
    red_mem[94] = 8'h00;
    red_mem[95] = 8'h00;
    red_mem[96] = 8'h00;
    red_mem[97] = 8'h00;
    red_mem[98] = 8'h00;
    red_mem[99] = 8'h00;
    red_mem[100] = 8'h00;
    red_mem[101] = 8'h00;
    red_mem[102] = 8'h00;
    red_mem[103] = 8'h00;
    red_mem[104] = 8'h00;
    red_mem[105] = 8'h00;
    red_mem[106] = 8'h00;
    red_mem[107] = 8'h00;
    red_mem[108] = 8'h00;
    red_mem[109] = 8'h00;
    red_mem[110] = 8'h00;
    red_mem[111] = 8'h00;
    red_mem[112] = 8'h00;
    red_mem[113] = 8'h00;
    red_mem[114] = 8'h00;
    red_mem[115] = 8'h00;
    red_mem[116] = 8'h00;
    red_mem[117] = 8'h00;
    red_mem[118] = 8'h00;
    red_mem[119] = 8'h00;
    red_mem[120] = 8'h00;
    red_mem[121] = 8'h00;
    red_mem[122] = 8'h00;
    red_mem[123] = 8'h00;
    red_mem[124] = 8'h00;
    red_mem[125] = 8'h00;
    red_mem[126] = 8'h00;
    red_mem[127] = 8'h00;
    red_mem[128] = 8'h00;
    red_mem[129] = 8'h00;
    red_mem[130] = 8'h00;
    red_mem[131] = 8'h00;
    red_mem[132] = 8'h00;
    red_mem[133] = 8'h00;
    red_mem[134] = 8'h00;
    red_mem[135] = 8'h00;
    red_mem[136] = 8'h00;
    red_mem[137] = 8'h00;
    red_mem[138] = 8'h00;
    red_mem[139] = 8'h00;
    red_mem[140] = 8'h00;
    red_mem[141] = 8'h00;
    red_mem[142] = 8'h00;
    red_mem[143] = 8'h00;
    red_mem[144] = 8'h00;
    red_mem[145] = 8'h00;
    red_mem[146] = 8'h00;
    red_mem[147] = 8'h00;
    red_mem[148] = 8'h00;
    red_mem[149] = 8'h00;
    red_mem[150] = 8'h00;
    red_mem[151] = 8'h00;
    red_mem[152] = 8'h00;
    red_mem[153] = 8'h00;
    red_mem[154] = 8'h00;
    red_mem[155] = 8'h00;
    red_mem[156] = 8'h00;
    red_mem[157] = 8'h00;
    red_mem[158] = 8'h00;
    red_mem[159] = 8'h00;
    red_mem[160] = 8'h00;
    red_mem[161] = 8'h00;
    red_mem[162] = 8'h00;
    red_mem[163] = 8'h00;
    red_mem[164] = 8'h00;
    red_mem[165] = 8'h00;
    red_mem[166] = 8'h00;
    red_mem[167] = 8'h00;
    red_mem[168] = 8'h00;
    red_mem[169] = 8'h00;
    red_mem[170] = 8'h00;
    red_mem[171] = 8'h00;
    red_mem[172] = 8'h00;
    red_mem[173] = 8'h00;
    red_mem[174] = 8'h00;
    red_mem[175] = 8'h00;
    red_mem[176] = 8'h00;
    red_mem[177] = 8'h00;
    red_mem[178] = 8'h00;
    red_mem[179] = 8'h00;
    red_mem[180] = 8'h00;
    red_mem[181] = 8'h00;
    red_mem[182] = 8'h00;
    red_mem[183] = 8'h00;
    red_mem[184] = 8'h00;
    red_mem[185] = 8'h00;
    red_mem[186] = 8'h00;
    red_mem[187] = 8'h00;
    red_mem[188] = 8'h00;
    red_mem[189] = 8'h00;
    red_mem[190] = 8'h00;
    red_mem[191] = 8'h00;
    red_mem[192] = 8'h00;
    red_mem[193] = 8'h00;
    red_mem[194] = 8'h00;
    red_mem[195] = 8'h00;
    red_mem[196] = 8'h00;
    red_mem[197] = 8'h00;
    red_mem[198] = 8'h00;
    red_mem[199] = 8'h00;
    red_mem[200] = 8'h00;
    red_mem[201] = 8'h00;
    red_mem[202] = 8'h00;
    red_mem[203] = 8'h00;
    red_mem[204] = 8'h00;
    red_mem[205] = 8'h00;
    red_mem[206] = 8'h00;
    red_mem[207] = 8'h00;
    red_mem[208] = 8'h00;
    red_mem[209] = 8'h00;
    red_mem[210] = 8'h00;
    red_mem[211] = 8'h00;
    red_mem[212] = 8'h00;
    red_mem[213] = 8'h00;
    red_mem[214] = 8'h00;
    red_mem[215] = 8'h00;
    red_mem[216] = 8'h00;
    red_mem[217] = 8'h00;
    red_mem[218] = 8'h00;
    red_mem[219] = 8'h00;
    red_mem[220] = 8'h00;
    red_mem[221] = 8'h00;
    red_mem[222] = 8'h00;
    red_mem[223] = 8'h00;
    red_mem[224] = 8'h00;
    red_mem[225] = 8'h00;
    red_mem[226] = 8'h00;
    red_mem[227] = 8'h00;
    red_mem[228] = 8'h00;
    red_mem[229] = 8'h00;
    red_mem[230] = 8'h00;
    red_mem[231] = 8'h00;
    red_mem[232] = 8'h00;
    red_mem[233] = 8'h00;
    red_mem[234] = 8'h00;
    red_mem[235] = 8'h00;
    red_mem[236] = 8'h00;
    red_mem[237] = 8'h00;
    red_mem[238] = 8'h00;
    red_mem[239] = 8'h00;
    red_mem[240] = 8'h00;
    red_mem[241] = 8'h00;
    red_mem[242] = 8'h00;
    red_mem[243] = 8'h00;
    red_mem[244] = 8'h00;
    red_mem[245] = 8'h00;
    red_mem[246] = 8'h00;
    red_mem[247] = 8'h00;
    red_mem[248] = 8'h00;
    red_mem[249] = 8'h00;
    red_mem[250] = 8'h00;
    red_mem[251] = 8'h00;
    red_mem[252] = 8'h00;
    red_mem[253] = 8'h00;
    red_mem[254] = 8'h00;
    red_mem[255] = 8'h00;
    red_mem[256] = 8'h00;
    red_mem[257] = 8'h00;
    red_mem[258] = 8'h00;
    red_mem[259] = 8'h00;
    red_mem[260] = 8'h00;
    red_mem[261] = 8'h00;
    red_mem[262] = 8'h00;
    red_mem[263] = 8'h00;
    red_mem[264] = 8'h00;
    red_mem[265] = 8'h00;
    red_mem[266] = 8'h00;
    red_mem[267] = 8'h00;
    red_mem[268] = 8'h00;
    red_mem[269] = 8'h00;
    red_mem[270] = 8'h00;
    red_mem[271] = 8'h00;
    red_mem[272] = 8'h00;
    red_mem[273] = 8'h00;
    red_mem[274] = 8'h00;
    red_mem[275] = 8'h00;
    red_mem[276] = 8'h00;
    red_mem[277] = 8'h00;
    red_mem[278] = 8'h00;
    red_mem[279] = 8'h00;
    red_mem[280] = 8'h00;
    red_mem[281] = 8'h00;
    red_mem[282] = 8'h00;
    red_mem[283] = 8'h00;
    red_mem[284] = 8'h00;
    red_mem[285] = 8'h00;
    red_mem[286] = 8'h00;
    red_mem[287] = 8'h00;
    red_mem[288] = 8'h00;
    red_mem[289] = 8'h00;
    red_mem[290] = 8'h00;
    red_mem[291] = 8'h00;
    red_mem[292] = 8'h00;
    red_mem[293] = 8'h00;
    red_mem[294] = 8'h00;
    red_mem[295] = 8'h00;
    red_mem[296] = 8'h00;
    red_mem[297] = 8'h00;
    red_mem[298] = 8'h00;
    red_mem[299] = 8'h00;
    red_mem[300] = 8'h00;
    red_mem[301] = 8'h00;
    red_mem[302] = 8'h00;
    red_mem[303] = 8'h00;
    red_mem[304] = 8'h00;
    red_mem[305] = 8'h00;
    red_mem[306] = 8'h00;
    red_mem[307] = 8'h00;
    red_mem[308] = 8'h00;
    red_mem[309] = 8'h00;
    red_mem[310] = 8'h00;
    red_mem[311] = 8'h00;
    red_mem[312] = 8'h00;
    red_mem[313] = 8'h00;
    red_mem[314] = 8'h00;
    red_mem[315] = 8'h00;
    red_mem[316] = 8'h00;
    red_mem[317] = 8'h00;
    red_mem[318] = 8'h00;
    red_mem[319] = 8'h00;
    red_mem[320] = 8'h00;
    red_mem[321] = 8'h00;
    red_mem[322] = 8'h00;
    red_mem[323] = 8'h00;
    red_mem[324] = 8'h00;
    red_mem[325] = 8'h00;
    red_mem[326] = 8'h00;
    red_mem[327] = 8'h00;
    red_mem[328] = 8'h00;
    red_mem[329] = 8'h00;
    red_mem[330] = 8'h00;
    red_mem[331] = 8'h00;
    red_mem[332] = 8'h00;
    red_mem[333] = 8'h00;
    red_mem[334] = 8'h00;
    red_mem[335] = 8'h00;
    red_mem[336] = 8'h00;
    red_mem[337] = 8'h00;
    red_mem[338] = 8'h00;
    red_mem[339] = 8'h00;
    red_mem[340] = 8'h00;
    red_mem[341] = 8'h00;
    red_mem[342] = 8'h00;
    red_mem[343] = 8'h00;
    red_mem[344] = 8'h00;
    red_mem[345] = 8'h00;
    red_mem[346] = 8'h00;
    red_mem[347] = 8'h00;
    red_mem[348] = 8'h00;
    red_mem[349] = 8'h00;
    red_mem[350] = 8'h00;
    red_mem[351] = 8'h00;
    red_mem[352] = 8'h00;
    red_mem[353] = 8'h00;
    red_mem[354] = 8'h00;
    red_mem[355] = 8'h00;
    red_mem[356] = 8'h00;
    red_mem[357] = 8'h00;
    red_mem[358] = 8'h00;
    red_mem[359] = 8'h00;
    red_mem[360] = 8'h00;
    red_mem[361] = 8'h00;
    red_mem[362] = 8'h00;
    red_mem[363] = 8'h00;
    red_mem[364] = 8'h00;
    red_mem[365] = 8'h00;
    red_mem[366] = 8'h00;
    red_mem[367] = 8'h00;
    red_mem[368] = 8'h00;
    red_mem[369] = 8'h00;
    red_mem[370] = 8'h00;
    red_mem[371] = 8'h00;
    red_mem[372] = 8'h00;
    red_mem[373] = 8'h00;
    red_mem[374] = 8'h00;
    red_mem[375] = 8'h00;
    red_mem[376] = 8'h00;
    red_mem[377] = 8'h00;
    red_mem[378] = 8'h00;
    red_mem[379] = 8'h00;
    red_mem[380] = 8'h00;
    red_mem[381] = 8'h00;
    red_mem[382] = 8'h00;
    red_mem[383] = 8'h00;
    red_mem[384] = 8'h00;
    red_mem[385] = 8'h00;
    red_mem[386] = 8'h00;
    red_mem[387] = 8'h00;
    red_mem[388] = 8'h00;
    red_mem[389] = 8'h00;
    red_mem[390] = 8'h00;
    red_mem[391] = 8'h00;
    red_mem[392] = 8'h00;
    red_mem[393] = 8'h00;
    red_mem[394] = 8'h00;
    red_mem[395] = 8'h00;
    red_mem[396] = 8'h00;
    red_mem[397] = 8'h00;
    red_mem[398] = 8'h00;
    red_mem[399] = 8'h00;
    red_mem[400] = 8'h00;
    red_mem[401] = 8'h00;
    red_mem[402] = 8'h00;
    red_mem[403] = 8'h00;
    red_mem[404] = 8'h00;
    red_mem[405] = 8'h00;
    red_mem[406] = 8'h00;
    red_mem[407] = 8'h00;
    red_mem[408] = 8'h00;
    red_mem[409] = 8'h00;
    red_mem[410] = 8'h00;
    red_mem[411] = 8'h00;
    red_mem[412] = 8'h00;
    red_mem[413] = 8'h00;
    red_mem[414] = 8'h00;
    red_mem[415] = 8'h00;
    red_mem[416] = 8'h00;
    red_mem[417] = 8'h00;
    red_mem[418] = 8'h00;
    red_mem[419] = 8'h00;
    red_mem[420] = 8'h00;
    red_mem[421] = 8'h00;
    red_mem[422] = 8'h00;
    red_mem[423] = 8'h00;
    red_mem[424] = 8'h00;
    red_mem[425] = 8'h00;
    red_mem[426] = 8'h00;
    red_mem[427] = 8'h00;
    red_mem[428] = 8'h00;
    red_mem[429] = 8'h00;
    red_mem[430] = 8'h00;
    red_mem[431] = 8'h00;
    red_mem[432] = 8'h00;
    red_mem[433] = 8'h00;
    red_mem[434] = 8'h00;
    red_mem[435] = 8'h00;
    red_mem[436] = 8'h00;
    red_mem[437] = 8'h00;
    red_mem[438] = 8'h00;
    red_mem[439] = 8'h00;
    red_mem[440] = 8'h00;
    red_mem[441] = 8'h00;
    red_mem[442] = 8'h00;
    red_mem[443] = 8'h00;
    red_mem[444] = 8'h00;
    red_mem[445] = 8'h00;
    red_mem[446] = 8'h00;
    red_mem[447] = 8'h00;
    red_mem[448] = 8'h00;
    red_mem[449] = 8'h00;
    red_mem[450] = 8'h00;
    red_mem[451] = 8'h00;
    red_mem[452] = 8'h00;
    red_mem[453] = 8'h00;
    red_mem[454] = 8'h00;
    red_mem[455] = 8'h00;
    red_mem[456] = 8'h00;
    red_mem[457] = 8'h00;
    red_mem[458] = 8'h00;
    red_mem[459] = 8'h00;
    red_mem[460] = 8'h00;
    red_mem[461] = 8'h00;
    red_mem[462] = 8'h00;
    red_mem[463] = 8'h00;
    red_mem[464] = 8'h00;
    red_mem[465] = 8'h00;
    red_mem[466] = 8'h00;
    red_mem[467] = 8'h00;
    red_mem[468] = 8'h00;
    red_mem[469] = 8'h00;
    red_mem[470] = 8'h00;
    red_mem[471] = 8'h00;
    red_mem[472] = 8'h00;
    red_mem[473] = 8'h00;
    red_mem[474] = 8'h00;
    red_mem[475] = 8'h00;
    red_mem[476] = 8'h00;
    red_mem[477] = 8'h00;
    red_mem[478] = 8'h00;
    red_mem[479] = 8'h00;
    red_mem[480] = 8'h00;
    red_mem[481] = 8'h00;
    red_mem[482] = 8'h00;
    red_mem[483] = 8'h00;
    red_mem[484] = 8'h00;
    red_mem[485] = 8'h00;
    red_mem[486] = 8'h00;
    red_mem[487] = 8'h00;
    red_mem[488] = 8'h00;
    red_mem[489] = 8'h00;
    red_mem[490] = 8'h00;
    red_mem[491] = 8'h00;
    red_mem[492] = 8'h00;
    red_mem[493] = 8'h00;
    red_mem[494] = 8'h00;
    red_mem[495] = 8'h00;
    red_mem[496] = 8'h00;
    red_mem[497] = 8'h00;
    red_mem[498] = 8'h00;
    red_mem[499] = 8'h00;
    red_mem[500] = 8'h00;
    red_mem[501] = 8'h00;
    red_mem[502] = 8'h00;
    red_mem[503] = 8'h00;
    red_mem[504] = 8'h00;
    red_mem[505] = 8'h00;
    red_mem[506] = 8'h00;
    red_mem[507] = 8'h00;
    red_mem[508] = 8'h00;
    red_mem[509] = 8'h00;
    red_mem[510] = 8'h00;
    red_mem[511] = 8'h00;
    red_mem[512] = 8'h00;
    red_mem[513] = 8'h00;
    red_mem[514] = 8'h00;
    red_mem[515] = 8'h00;
    red_mem[516] = 8'h00;
    red_mem[517] = 8'h00;
    red_mem[518] = 8'h00;
    red_mem[519] = 8'h00;
    red_mem[520] = 8'h00;
    red_mem[521] = 8'h00;
    red_mem[522] = 8'h00;
    red_mem[523] = 8'h00;
    red_mem[524] = 8'h00;
    red_mem[525] = 8'h00;
    red_mem[526] = 8'h00;
    red_mem[527] = 8'h00;
    red_mem[528] = 8'h00;
    red_mem[529] = 8'h00;
    red_mem[530] = 8'h00;
    red_mem[531] = 8'h00;
    red_mem[532] = 8'h00;
    red_mem[533] = 8'h00;
    red_mem[534] = 8'h00;
    red_mem[535] = 8'h00;
    red_mem[536] = 8'h00;
    red_mem[537] = 8'h00;
    red_mem[538] = 8'h00;
    red_mem[539] = 8'h00;
    red_mem[540] = 8'h00;
    red_mem[541] = 8'h00;
    red_mem[542] = 8'h00;
    red_mem[543] = 8'h00;
    red_mem[544] = 8'h00;
    red_mem[545] = 8'h00;
    red_mem[546] = 8'h00;
    red_mem[547] = 8'h00;
    red_mem[548] = 8'h00;
    red_mem[549] = 8'h00;
    red_mem[550] = 8'h00;
    red_mem[551] = 8'h00;
    red_mem[552] = 8'h00;
    red_mem[553] = 8'h00;
    red_mem[554] = 8'h00;
    red_mem[555] = 8'h00;
    red_mem[556] = 8'h00;
    red_mem[557] = 8'h00;
    red_mem[558] = 8'h00;
    red_mem[559] = 8'h00;
    red_mem[560] = 8'h00;
    red_mem[561] = 8'h00;
    red_mem[562] = 8'h00;
    red_mem[563] = 8'h00;
    red_mem[564] = 8'h00;
    red_mem[565] = 8'h00;
    red_mem[566] = 8'h00;
    red_mem[567] = 8'h00;
    red_mem[568] = 8'h00;
    red_mem[569] = 8'h00;
    red_mem[570] = 8'h00;
    red_mem[571] = 8'h00;
    red_mem[572] = 8'h00;
    red_mem[573] = 8'h00;
    red_mem[574] = 8'h00;
    red_mem[575] = 8'h00;
    red_mem[576] = 8'h00;
    red_mem[577] = 8'h00;
    red_mem[578] = 8'h00;
    red_mem[579] = 8'h00;
    red_mem[580] = 8'h00;
    red_mem[581] = 8'h00;
    red_mem[582] = 8'h00;
    red_mem[583] = 8'h00;
    red_mem[584] = 8'h00;
    red_mem[585] = 8'h00;
    red_mem[586] = 8'h00;
    red_mem[587] = 8'h00;
    red_mem[588] = 8'h00;
    red_mem[589] = 8'h00;
    red_mem[590] = 8'h00;
    red_mem[591] = 8'h00;
    red_mem[592] = 8'h00;
    red_mem[593] = 8'h00;
    red_mem[594] = 8'h00;
    red_mem[595] = 8'h00;
    red_mem[596] = 8'h00;
    red_mem[597] = 8'h00;
    red_mem[598] = 8'he0;
    red_mem[599] = 8'h00;
    red_mem[600] = 8'h00;
    red_mem[601] = 8'he0;
    red_mem[602] = 8'h3b;
    red_mem[603] = 8'h00;
    red_mem[604] = 8'h00;
    red_mem[605] = 8'h00;
    red_mem[606] = 8'h00;
    red_mem[607] = 8'h00;
    red_mem[608] = 8'h00;
    red_mem[609] = 8'h00;
    red_mem[610] = 8'h00;
    red_mem[611] = 8'h00;
    red_mem[612] = 8'h00;
    red_mem[613] = 8'h00;
    red_mem[614] = 8'hf8;
    red_mem[615] = 8'h00;
    red_mem[616] = 8'h00;
    red_mem[617] = 8'hfe;
    red_mem[618] = 8'hff;
    red_mem[619] = 8'h03;
    red_mem[620] = 8'h00;
    red_mem[621] = 8'h00;
    red_mem[622] = 8'h00;
    red_mem[623] = 8'h00;
    red_mem[624] = 8'h00;
    red_mem[625] = 8'h00;
    red_mem[626] = 8'h00;
    red_mem[627] = 8'h00;
    red_mem[628] = 8'h00;
    red_mem[629] = 8'h00;
    red_mem[630] = 8'hfc;
    red_mem[631] = 8'h00;
    red_mem[632] = 8'h00;
    red_mem[633] = 8'hff;
    red_mem[634] = 8'hff;
    red_mem[635] = 8'h0f;
    red_mem[636] = 8'h00;
    red_mem[637] = 8'h00;
    red_mem[638] = 8'h00;
    red_mem[639] = 8'h00;
    red_mem[640] = 8'h00;
    red_mem[641] = 8'h00;
    red_mem[642] = 8'h00;
    red_mem[643] = 8'h00;
    red_mem[644] = 8'h00;
    red_mem[645] = 8'h00;
    red_mem[646] = 8'h7e;
    red_mem[647] = 8'h00;
    red_mem[648] = 8'hc0;
    red_mem[649] = 8'hff;
    red_mem[650] = 8'hff;
    red_mem[651] = 8'h0f;
    red_mem[652] = 8'h00;
    red_mem[653] = 8'h00;
    red_mem[654] = 8'h00;
    red_mem[655] = 8'h00;
    red_mem[656] = 8'h00;
    red_mem[657] = 8'h00;
    red_mem[658] = 8'h00;
    red_mem[659] = 8'h00;
    red_mem[660] = 8'h00;
    red_mem[661] = 8'h00;
    red_mem[662] = 8'hff;
    red_mem[663] = 8'h00;
    red_mem[664] = 8'hc0;
    red_mem[665] = 8'h0f;
    red_mem[666] = 8'hfe;
    red_mem[667] = 8'h1f;
    red_mem[668] = 8'h00;
    red_mem[669] = 8'h00;
    red_mem[670] = 8'h00;
    red_mem[671] = 8'h00;
    red_mem[672] = 8'h00;
    red_mem[673] = 8'h00;
    red_mem[674] = 8'h00;
    red_mem[675] = 8'h00;
    red_mem[676] = 8'h00;
    red_mem[677] = 8'h00;
    red_mem[678] = 8'hff;
    red_mem[679] = 8'h00;
    red_mem[680] = 8'hf8;
    red_mem[681] = 8'h07;
    red_mem[682] = 8'hf8;
    red_mem[683] = 8'h1f;
    red_mem[684] = 8'h00;
    red_mem[685] = 8'h00;
    red_mem[686] = 8'h00;
    red_mem[687] = 8'h00;
    red_mem[688] = 8'h00;
    red_mem[689] = 8'h00;
    red_mem[690] = 8'h00;
    red_mem[691] = 8'h00;
    red_mem[692] = 8'h00;
    red_mem[693] = 8'hc0;
    red_mem[694] = 8'h7f;
    red_mem[695] = 8'h00;
    red_mem[696] = 8'hf8;
    red_mem[697] = 8'h03;
    red_mem[698] = 8'hc0;
    red_mem[699] = 8'h1f;
    red_mem[700] = 8'h00;
    red_mem[701] = 8'h00;
    red_mem[702] = 8'h00;
    red_mem[703] = 8'h00;
    red_mem[704] = 8'h00;
    red_mem[705] = 8'h00;
    red_mem[706] = 8'h00;
    red_mem[707] = 8'h00;
    red_mem[708] = 8'h00;
    red_mem[709] = 8'hc0;
    red_mem[710] = 8'h7f;
    red_mem[711] = 8'h00;
    red_mem[712] = 8'hfc;
    red_mem[713] = 8'h01;
    red_mem[714] = 8'h80;
    red_mem[715] = 8'h3f;
    red_mem[716] = 8'h00;
    red_mem[717] = 8'h00;
    red_mem[718] = 8'h00;
    red_mem[719] = 8'h00;
    red_mem[720] = 8'h00;
    red_mem[721] = 8'h00;
    red_mem[722] = 8'h00;
    red_mem[723] = 8'h00;
    red_mem[724] = 8'h00;
    red_mem[725] = 8'hf0;
    red_mem[726] = 8'h3f;
    red_mem[727] = 8'h00;
    red_mem[728] = 8'hfc;
    red_mem[729] = 8'h00;
    red_mem[730] = 8'h80;
    red_mem[731] = 8'h7f;
    red_mem[732] = 8'h00;
    red_mem[733] = 8'h00;
    red_mem[734] = 8'h00;
    red_mem[735] = 8'h00;
    red_mem[736] = 8'h00;
    red_mem[737] = 8'h00;
    red_mem[738] = 8'h00;
    red_mem[739] = 8'h00;
    red_mem[740] = 8'h00;
    red_mem[741] = 8'hf0;
    red_mem[742] = 8'h7f;
    red_mem[743] = 8'h00;
    red_mem[744] = 8'hfe;
    red_mem[745] = 8'h00;
    red_mem[746] = 8'h00;
    red_mem[747] = 8'h7f;
    red_mem[748] = 8'h00;
    red_mem[749] = 8'h00;
    red_mem[750] = 8'h00;
    red_mem[751] = 8'h00;
    red_mem[752] = 8'h00;
    red_mem[753] = 8'h00;
    red_mem[754] = 8'h00;
    red_mem[755] = 8'h00;
    red_mem[756] = 8'h00;
    red_mem[757] = 8'hf0;
    red_mem[758] = 8'h3f;
    red_mem[759] = 8'h00;
    red_mem[760] = 8'hfc;
    red_mem[761] = 8'h00;
    red_mem[762] = 8'h00;
    red_mem[763] = 8'hff;
    red_mem[764] = 8'h00;
    red_mem[765] = 8'h00;
    red_mem[766] = 8'h00;
    red_mem[767] = 8'h00;
    red_mem[768] = 8'h00;
    red_mem[769] = 8'h00;
    red_mem[770] = 8'h00;
    red_mem[771] = 8'h00;
    red_mem[772] = 8'h00;
    red_mem[773] = 8'hfe;
    red_mem[774] = 8'h1f;
    red_mem[775] = 8'h00;
    red_mem[776] = 8'hfe;
    red_mem[777] = 8'h00;
    red_mem[778] = 8'h80;
    red_mem[779] = 8'hff;
    red_mem[780] = 8'h00;
    red_mem[781] = 8'h00;
    red_mem[782] = 8'h00;
    red_mem[783] = 8'h00;
    red_mem[784] = 8'h00;
    red_mem[785] = 8'h00;
    red_mem[786] = 8'h00;
    red_mem[787] = 8'h00;
    red_mem[788] = 8'h00;
    red_mem[789] = 8'h9e;
    red_mem[790] = 8'h3f;
    red_mem[791] = 8'h00;
    red_mem[792] = 8'hfe;
    red_mem[793] = 8'h01;
    red_mem[794] = 8'h80;
    red_mem[795] = 8'hff;
    red_mem[796] = 8'h00;
    red_mem[797] = 8'h00;
    red_mem[798] = 8'h00;
    red_mem[799] = 8'h00;
    red_mem[800] = 8'h00;
    red_mem[801] = 8'h00;
    red_mem[802] = 8'h00;
    red_mem[803] = 8'h00;
    red_mem[804] = 8'hc0;
    red_mem[805] = 8'h8f;
    red_mem[806] = 8'h3f;
    red_mem[807] = 8'h00;
    red_mem[808] = 8'hff;
    red_mem[809] = 8'h07;
    red_mem[810] = 8'h00;
    red_mem[811] = 8'hff;
    red_mem[812] = 8'h00;
    red_mem[813] = 8'h00;
    red_mem[814] = 8'h00;
    red_mem[815] = 8'h00;
    red_mem[816] = 8'h00;
    red_mem[817] = 8'h00;
    red_mem[818] = 8'h00;
    red_mem[819] = 8'h00;
    red_mem[820] = 8'hc0;
    red_mem[821] = 8'h8f;
    red_mem[822] = 8'h1f;
    red_mem[823] = 8'h00;
    red_mem[824] = 8'hfb;
    red_mem[825] = 8'h07;
    red_mem[826] = 8'hc0;
    red_mem[827] = 8'hff;
    red_mem[828] = 8'h00;
    red_mem[829] = 8'h00;
    red_mem[830] = 8'h00;
    red_mem[831] = 8'h00;
    red_mem[832] = 8'h00;
    red_mem[833] = 8'h00;
    red_mem[834] = 8'h00;
    red_mem[835] = 8'h00;
    red_mem[836] = 8'hc0;
    red_mem[837] = 8'hc7;
    red_mem[838] = 8'h1d;
    red_mem[839] = 8'h00;
    red_mem[840] = 8'hff;
    red_mem[841] = 8'h0f;
    red_mem[842] = 8'hc0;
    red_mem[843] = 8'hff;
    red_mem[844] = 8'h00;
    red_mem[845] = 8'h00;
    red_mem[846] = 8'h00;
    red_mem[847] = 8'h00;
    red_mem[848] = 8'h00;
    red_mem[849] = 8'h00;
    red_mem[850] = 8'h00;
    red_mem[851] = 8'h00;
    red_mem[852] = 8'hc0;
    red_mem[853] = 8'hc3;
    red_mem[854] = 8'h1f;
    red_mem[855] = 8'h00;
    red_mem[856] = 8'hff;
    red_mem[857] = 8'h07;
    red_mem[858] = 8'hc0;
    red_mem[859] = 8'h7f;
    red_mem[860] = 8'h00;
    red_mem[861] = 8'h00;
    red_mem[862] = 8'h00;
    red_mem[863] = 8'h00;
    red_mem[864] = 8'h00;
    red_mem[865] = 8'h00;
    red_mem[866] = 8'h00;
    red_mem[867] = 8'h00;
    red_mem[868] = 8'hc0;
    red_mem[869] = 8'hc1;
    red_mem[870] = 8'h1f;
    red_mem[871] = 8'h00;
    red_mem[872] = 8'hff;
    red_mem[873] = 8'h05;
    red_mem[874] = 8'hc0;
    red_mem[875] = 8'h7f;
    red_mem[876] = 8'h00;
    red_mem[877] = 8'h00;
    red_mem[878] = 8'h00;
    red_mem[879] = 8'h00;
    red_mem[880] = 8'h00;
    red_mem[881] = 8'h00;
    red_mem[882] = 8'h00;
    red_mem[883] = 8'h00;
    red_mem[884] = 8'h00;
    red_mem[885] = 8'he0;
    red_mem[886] = 8'h0f;
    red_mem[887] = 8'h00;
    red_mem[888] = 8'hff;
    red_mem[889] = 8'h07;
    red_mem[890] = 8'he0;
    red_mem[891] = 8'h7f;
    red_mem[892] = 8'h00;
    red_mem[893] = 8'h00;
    red_mem[894] = 8'h00;
    red_mem[895] = 8'h00;
    red_mem[896] = 8'h00;
    red_mem[897] = 8'h00;
    red_mem[898] = 8'h00;
    red_mem[899] = 8'h00;
    red_mem[900] = 8'h00;
    red_mem[901] = 8'he0;
    red_mem[902] = 8'h0f;
    red_mem[903] = 8'h00;
    red_mem[904] = 8'hfc;
    red_mem[905] = 8'h07;
    red_mem[906] = 8'he0;
    red_mem[907] = 8'h7f;
    red_mem[908] = 8'h00;
    red_mem[909] = 8'h00;
    red_mem[910] = 8'h00;
    red_mem[911] = 8'h00;
    red_mem[912] = 8'h00;
    red_mem[913] = 8'h00;
    red_mem[914] = 8'h00;
    red_mem[915] = 8'h00;
    red_mem[916] = 8'h00;
    red_mem[917] = 8'he0;
    red_mem[918] = 8'h1f;
    red_mem[919] = 8'h00;
    red_mem[920] = 8'hfc;
    red_mem[921] = 8'h01;
    red_mem[922] = 8'hf0;
    red_mem[923] = 8'h0f;
    red_mem[924] = 8'h00;
    red_mem[925] = 8'h00;
    red_mem[926] = 8'h00;
    red_mem[927] = 8'h00;
    red_mem[928] = 8'h00;
    red_mem[929] = 8'h00;
    red_mem[930] = 8'h00;
    red_mem[931] = 8'h00;
    red_mem[932] = 8'h00;
    red_mem[933] = 8'hf0;
    red_mem[934] = 8'h0f;
    red_mem[935] = 8'h00;
    red_mem[936] = 8'h60;
    red_mem[937] = 8'h00;
    red_mem[938] = 8'hf8;
    red_mem[939] = 8'h0f;
    red_mem[940] = 8'h00;
    red_mem[941] = 8'h00;
    red_mem[942] = 8'h00;
    red_mem[943] = 8'h00;
    red_mem[944] = 8'h00;
    red_mem[945] = 8'h00;
    red_mem[946] = 8'h00;
    red_mem[947] = 8'h00;
    red_mem[948] = 8'h00;
    red_mem[949] = 8'hf0;
    red_mem[950] = 8'h0f;
    red_mem[951] = 8'h00;
    red_mem[952] = 8'h00;
    red_mem[953] = 8'h00;
    red_mem[954] = 8'hff;
    red_mem[955] = 8'h07;
    red_mem[956] = 8'h00;
    red_mem[957] = 8'h00;
    red_mem[958] = 8'h00;
    red_mem[959] = 8'h00;
    red_mem[960] = 8'h00;
    red_mem[961] = 8'h00;
    red_mem[962] = 8'h00;
    red_mem[963] = 8'h00;
    red_mem[964] = 8'h00;
    red_mem[965] = 8'he0;
    red_mem[966] = 8'h07;
    red_mem[967] = 8'h00;
    red_mem[968] = 8'h00;
    red_mem[969] = 8'h80;
    red_mem[970] = 8'hff;
    red_mem[971] = 8'h03;
    red_mem[972] = 8'h00;
    red_mem[973] = 8'h00;
    red_mem[974] = 8'h00;
    red_mem[975] = 8'h00;
    red_mem[976] = 8'h00;
    red_mem[977] = 8'h00;
    red_mem[978] = 8'h00;
    red_mem[979] = 8'h00;
    red_mem[980] = 8'h00;
    red_mem[981] = 8'hf0;
    red_mem[982] = 8'h07;
    red_mem[983] = 8'h00;
    red_mem[984] = 8'h00;
    red_mem[985] = 8'h80;
    red_mem[986] = 8'hff;
    red_mem[987] = 8'h00;
    red_mem[988] = 8'h00;
    red_mem[989] = 8'h00;
    red_mem[990] = 8'h00;
    red_mem[991] = 8'h00;
    red_mem[992] = 8'h00;
    red_mem[993] = 8'h00;
    red_mem[994] = 8'h00;
    red_mem[995] = 8'h00;
    red_mem[996] = 8'h00;
    red_mem[997] = 8'hf0;
    red_mem[998] = 8'h07;
    red_mem[999] = 8'h00;
    red_mem[1000] = 8'h00;
    red_mem[1001] = 8'h80;
    red_mem[1002] = 8'hff;
    red_mem[1003] = 8'h00;
    red_mem[1004] = 8'h00;
    red_mem[1005] = 8'h00;
    red_mem[1006] = 8'h00;
    red_mem[1007] = 8'h00;
    red_mem[1008] = 8'h00;
    red_mem[1009] = 8'h00;
    red_mem[1010] = 8'h00;
    red_mem[1011] = 8'h00;
    red_mem[1012] = 8'h00;
    red_mem[1013] = 8'hf0;
    red_mem[1014] = 8'h07;
    red_mem[1015] = 8'h00;
    red_mem[1016] = 8'h00;
    red_mem[1017] = 8'he0;
    red_mem[1018] = 8'h1f;
    red_mem[1019] = 8'h00;
    red_mem[1020] = 8'h00;
    red_mem[1021] = 8'h00;
    red_mem[1022] = 8'h00;
    red_mem[1023] = 8'h00;
    red_mem[1024] = 8'h00;
    red_mem[1025] = 8'h00;
    red_mem[1026] = 8'h00;
    red_mem[1027] = 8'h00;
    red_mem[1028] = 8'h00;
    red_mem[1029] = 8'hf8;
    red_mem[1030] = 8'h07;
    red_mem[1031] = 8'h00;
    red_mem[1032] = 8'h00;
    red_mem[1033] = 8'hf8;
    red_mem[1034] = 8'h0f;
    red_mem[1035] = 8'h00;
    red_mem[1036] = 8'h00;
    red_mem[1037] = 8'h00;
    red_mem[1038] = 8'h00;
    red_mem[1039] = 8'h00;
    red_mem[1040] = 8'h00;
    red_mem[1041] = 8'h00;
    red_mem[1042] = 8'h00;
    red_mem[1043] = 8'h00;
    red_mem[1044] = 8'h00;
    red_mem[1045] = 8'hf8;
    red_mem[1046] = 8'h07;
    red_mem[1047] = 8'h00;
    red_mem[1048] = 8'h00;
    red_mem[1049] = 8'hfc;
    red_mem[1050] = 8'h01;
    red_mem[1051] = 8'h00;
    red_mem[1052] = 8'h00;
    red_mem[1053] = 8'h00;
    red_mem[1054] = 8'h00;
    red_mem[1055] = 8'h00;
    red_mem[1056] = 8'h00;
    red_mem[1057] = 8'h00;
    red_mem[1058] = 8'h00;
    red_mem[1059] = 8'h00;
    red_mem[1060] = 8'h00;
    red_mem[1061] = 8'hf8;
    red_mem[1062] = 8'h03;
    red_mem[1063] = 8'h00;
    red_mem[1064] = 8'h00;
    red_mem[1065] = 8'hbe;
    red_mem[1066] = 8'h00;
    red_mem[1067] = 8'h00;
    red_mem[1068] = 8'h00;
    red_mem[1069] = 8'h00;
    red_mem[1070] = 8'h00;
    red_mem[1071] = 8'h00;
    red_mem[1072] = 8'h00;
    red_mem[1073] = 8'h00;
    red_mem[1074] = 8'h00;
    red_mem[1075] = 8'h00;
    red_mem[1076] = 8'h00;
    red_mem[1077] = 8'hfc;
    red_mem[1078] = 8'h01;
    red_mem[1079] = 8'h00;
    red_mem[1080] = 8'h80;
    red_mem[1081] = 8'h1f;
    red_mem[1082] = 8'h00;
    red_mem[1083] = 8'h00;
    red_mem[1084] = 8'h00;
    red_mem[1085] = 8'h00;
    red_mem[1086] = 8'h00;
    red_mem[1087] = 8'h00;
    red_mem[1088] = 8'h00;
    red_mem[1089] = 8'h00;
    red_mem[1090] = 8'h00;
    red_mem[1091] = 8'h00;
    red_mem[1092] = 8'h00;
    red_mem[1093] = 8'hfc;
    red_mem[1094] = 8'h01;
    red_mem[1095] = 8'h00;
    red_mem[1096] = 8'hc0;
    red_mem[1097] = 8'h1f;
    red_mem[1098] = 8'h00;
    red_mem[1099] = 8'h00;
    red_mem[1100] = 8'h00;
    red_mem[1101] = 8'h00;
    red_mem[1102] = 8'h00;
    red_mem[1103] = 8'h00;
    red_mem[1104] = 8'h00;
    red_mem[1105] = 8'h00;
    red_mem[1106] = 8'h00;
    red_mem[1107] = 8'h00;
    red_mem[1108] = 8'h00;
    red_mem[1109] = 8'hfc;
    red_mem[1110] = 8'h01;
    red_mem[1111] = 8'h00;
    red_mem[1112] = 8'he0;
    red_mem[1113] = 8'h03;
    red_mem[1114] = 8'h00;
    red_mem[1115] = 8'h00;
    red_mem[1116] = 8'h00;
    red_mem[1117] = 8'h00;
    red_mem[1118] = 8'h00;
    red_mem[1119] = 8'h00;
    red_mem[1120] = 8'h00;
    red_mem[1121] = 8'h00;
    red_mem[1122] = 8'h00;
    red_mem[1123] = 8'h00;
    red_mem[1124] = 8'h00;
    red_mem[1125] = 8'hfc;
    red_mem[1126] = 8'h00;
    red_mem[1127] = 8'h00;
    red_mem[1128] = 8'hf8;
    red_mem[1129] = 8'h03;
    red_mem[1130] = 8'h00;
    red_mem[1131] = 8'h00;
    red_mem[1132] = 8'h00;
    red_mem[1133] = 8'h00;
    red_mem[1134] = 8'h00;
    red_mem[1135] = 8'h00;
    red_mem[1136] = 8'h00;
    red_mem[1137] = 8'h00;
    red_mem[1138] = 8'h00;
    red_mem[1139] = 8'h00;
    red_mem[1140] = 8'h00;
    red_mem[1141] = 8'hfc;
    red_mem[1142] = 8'h01;
    red_mem[1143] = 8'h00;
    red_mem[1144] = 8'h78;
    red_mem[1145] = 8'h00;
    red_mem[1146] = 8'h00;
    red_mem[1147] = 8'h00;
    red_mem[1148] = 8'h00;
    red_mem[1149] = 8'h00;
    red_mem[1150] = 8'h00;
    red_mem[1151] = 8'h00;
    red_mem[1152] = 8'h00;
    red_mem[1153] = 8'h00;
    red_mem[1154] = 8'h00;
    red_mem[1155] = 8'h00;
    red_mem[1156] = 8'h00;
    red_mem[1157] = 8'hfe;
    red_mem[1158] = 8'h01;
    red_mem[1159] = 8'h00;
    red_mem[1160] = 8'h7f;
    red_mem[1161] = 8'h00;
    red_mem[1162] = 8'h00;
    red_mem[1163] = 8'h00;
    red_mem[1164] = 8'h00;
    red_mem[1165] = 8'h00;
    red_mem[1166] = 8'h00;
    red_mem[1167] = 8'h00;
    red_mem[1168] = 8'h00;
    red_mem[1169] = 8'h00;
    red_mem[1170] = 8'h00;
    red_mem[1171] = 8'h00;
    red_mem[1172] = 8'h00;
    red_mem[1173] = 8'hfc;
    red_mem[1174] = 8'h01;
    red_mem[1175] = 8'h80;
    red_mem[1176] = 8'hff;
    red_mem[1177] = 8'h02;
    red_mem[1178] = 8'h00;
    red_mem[1179] = 8'h00;
    red_mem[1180] = 8'h00;
    red_mem[1181] = 8'h00;
    red_mem[1182] = 8'h00;
    red_mem[1183] = 8'h00;
    red_mem[1184] = 8'h00;
    red_mem[1185] = 8'h00;
    red_mem[1186] = 8'h00;
    red_mem[1187] = 8'h00;
    red_mem[1188] = 8'h00;
    red_mem[1189] = 8'hfc;
    red_mem[1190] = 8'h01;
    red_mem[1191] = 8'h80;
    red_mem[1192] = 8'hff;
    red_mem[1193] = 8'h07;
    red_mem[1194] = 8'h00;
    red_mem[1195] = 8'h18;
    red_mem[1196] = 8'h00;
    red_mem[1197] = 8'h00;
    red_mem[1198] = 8'h00;
    red_mem[1199] = 8'h00;
    red_mem[1200] = 8'h00;
    red_mem[1201] = 8'h00;
    red_mem[1202] = 8'h00;
    red_mem[1203] = 8'h00;
    red_mem[1204] = 8'h00;
    red_mem[1205] = 8'hf8;
    red_mem[1206] = 8'h00;
    red_mem[1207] = 8'h80;
    red_mem[1208] = 8'hff;
    red_mem[1209] = 8'h7f;
    red_mem[1210] = 8'h00;
    red_mem[1211] = 8'h1c;
    red_mem[1212] = 8'h00;
    red_mem[1213] = 8'h00;
    red_mem[1214] = 8'h00;
    red_mem[1215] = 8'h00;
    red_mem[1216] = 8'h00;
    red_mem[1217] = 8'h00;
    red_mem[1218] = 8'h00;
    red_mem[1219] = 8'h00;
    red_mem[1220] = 8'h00;
    red_mem[1221] = 8'hfe;
    red_mem[1222] = 8'h00;
    red_mem[1223] = 8'hf0;
    red_mem[1224] = 8'hff;
    red_mem[1225] = 8'hff;
    red_mem[1226] = 8'h07;
    red_mem[1227] = 8'h0e;
    red_mem[1228] = 8'h00;
    red_mem[1229] = 8'h00;
    red_mem[1230] = 8'h00;
    red_mem[1231] = 8'h00;
    red_mem[1232] = 8'h00;
    red_mem[1233] = 8'h00;
    red_mem[1234] = 8'h00;
    red_mem[1235] = 8'h00;
    red_mem[1236] = 8'h00;
    red_mem[1237] = 8'h6f;
    red_mem[1238] = 8'h00;
    red_mem[1239] = 8'hf8;
    red_mem[1240] = 8'hff;
    red_mem[1241] = 8'hff;
    red_mem[1242] = 8'he7;
    red_mem[1243] = 8'h0f;
    red_mem[1244] = 8'h00;
    red_mem[1245] = 8'h00;
    red_mem[1246] = 8'h00;
    red_mem[1247] = 8'h00;
    red_mem[1248] = 8'h00;
    red_mem[1249] = 8'h00;
    red_mem[1250] = 8'h00;
    red_mem[1251] = 8'h00;
    red_mem[1252] = 8'h00;
    red_mem[1253] = 8'h7f;
    red_mem[1254] = 8'h00;
    red_mem[1255] = 8'hf8;
    red_mem[1256] = 8'hff;
    red_mem[1257] = 8'hff;
    red_mem[1258] = 8'hef;
    red_mem[1259] = 8'h07;
    red_mem[1260] = 8'h00;
    red_mem[1261] = 8'h00;
    red_mem[1262] = 8'h00;
    red_mem[1263] = 8'h00;
    red_mem[1264] = 8'h00;
    red_mem[1265] = 8'h00;
    red_mem[1266] = 8'h00;
    red_mem[1267] = 8'h00;
    red_mem[1268] = 8'h00;
    red_mem[1269] = 8'h7f;
    red_mem[1270] = 8'h00;
    red_mem[1271] = 8'hf8;
    red_mem[1272] = 8'hff;
    red_mem[1273] = 8'hff;
    red_mem[1274] = 8'hff;
    red_mem[1275] = 8'h07;
    red_mem[1276] = 8'h00;
    red_mem[1277] = 8'h00;
    red_mem[1278] = 8'h00;
    red_mem[1279] = 8'h00;
    red_mem[1280] = 8'h00;
    red_mem[1281] = 8'h00;
    red_mem[1282] = 8'h00;
    red_mem[1283] = 8'h00;
    red_mem[1284] = 8'h00;
    red_mem[1285] = 8'hff;
    red_mem[1286] = 8'h00;
    red_mem[1287] = 8'hf8;
    red_mem[1288] = 8'he6;
    red_mem[1289] = 8'hbf;
    red_mem[1290] = 8'hff;
    red_mem[1291] = 8'h03;
    red_mem[1292] = 8'h00;
    red_mem[1293] = 8'h00;
    red_mem[1294] = 8'h00;
    red_mem[1295] = 8'h00;
    red_mem[1296] = 8'h00;
    red_mem[1297] = 8'h00;
    red_mem[1298] = 8'h00;
    red_mem[1299] = 8'h00;
    red_mem[1300] = 8'hc8;
    red_mem[1301] = 8'hff;
    red_mem[1302] = 8'h07;
    red_mem[1303] = 8'h7f;
    red_mem[1304] = 8'h00;
    red_mem[1305] = 8'hfe;
    red_mem[1306] = 8'hff;
    red_mem[1307] = 8'h03;
    red_mem[1308] = 8'h00;
    red_mem[1309] = 8'h00;
    red_mem[1310] = 8'h00;
    red_mem[1311] = 8'h00;
    red_mem[1312] = 8'h00;
    red_mem[1313] = 8'h00;
    red_mem[1314] = 8'h00;
    red_mem[1315] = 8'h00;
    red_mem[1316] = 8'hfc;
    red_mem[1317] = 8'hff;
    red_mem[1318] = 8'h0f;
    red_mem[1319] = 8'h0f;
    red_mem[1320] = 8'h00;
    red_mem[1321] = 8'hfe;
    red_mem[1322] = 8'hff;
    red_mem[1323] = 8'h01;
    red_mem[1324] = 8'h00;
    red_mem[1325] = 8'h00;
    red_mem[1326] = 8'h00;
    red_mem[1327] = 8'h00;
    red_mem[1328] = 8'h00;
    red_mem[1329] = 8'h00;
    red_mem[1330] = 8'h00;
    red_mem[1331] = 8'h00;
    red_mem[1332] = 8'hfc;
    red_mem[1333] = 8'hff;
    red_mem[1334] = 8'h0f;
    red_mem[1335] = 8'h0f;
    red_mem[1336] = 8'h00;
    red_mem[1337] = 8'hf0;
    red_mem[1338] = 8'h3f;
    red_mem[1339] = 8'h00;
    red_mem[1340] = 8'h00;
    red_mem[1341] = 8'h00;
    red_mem[1342] = 8'h00;
    red_mem[1343] = 8'h00;
    red_mem[1344] = 8'h00;
    red_mem[1345] = 8'h00;
    red_mem[1346] = 8'h00;
    red_mem[1347] = 8'h00;
    red_mem[1348] = 8'hdc;
    red_mem[1349] = 8'h79;
    red_mem[1350] = 8'h0f;
    red_mem[1351] = 8'h06;
    red_mem[1352] = 8'h00;
    red_mem[1353] = 8'h00;
    red_mem[1354] = 8'h07;
    red_mem[1355] = 8'h00;
    red_mem[1356] = 8'h00;
    red_mem[1357] = 8'h00;
    red_mem[1358] = 8'h00;
    red_mem[1359] = 8'h00;
    red_mem[1360] = 8'h00;
    red_mem[1361] = 8'h00;
    red_mem[1362] = 8'h00;
    red_mem[1363] = 8'h00;
    red_mem[1364] = 8'h00;
    red_mem[1365] = 8'h00;
    red_mem[1366] = 8'h00;
    red_mem[1367] = 8'h00;
    red_mem[1368] = 8'h00;
    red_mem[1369] = 8'h00;
    red_mem[1370] = 8'h00;
    red_mem[1371] = 8'h00;
    red_mem[1372] = 8'h00;
    red_mem[1373] = 8'h00;
    red_mem[1374] = 8'h00;
    red_mem[1375] = 8'h00;
    red_mem[1376] = 8'h00;
    red_mem[1377] = 8'h00;
    red_mem[1378] = 8'h00;
    red_mem[1379] = 8'h00;
    red_mem[1380] = 8'h00;
    red_mem[1381] = 8'h00;
    red_mem[1382] = 8'h00;
    red_mem[1383] = 8'h00;
    red_mem[1384] = 8'h00;
    red_mem[1385] = 8'h00;
    red_mem[1386] = 8'h00;
    red_mem[1387] = 8'h00;
    red_mem[1388] = 8'h00;
    red_mem[1389] = 8'h00;
    red_mem[1390] = 8'h00;
    red_mem[1391] = 8'h00;
    red_mem[1392] = 8'h00;
    red_mem[1393] = 8'h00;
    red_mem[1394] = 8'h00;
    red_mem[1395] = 8'h00;
    red_mem[1396] = 8'h00;
    red_mem[1397] = 8'h00;
    red_mem[1398] = 8'h00;
    red_mem[1399] = 8'h00;
    red_mem[1400] = 8'h00;
    red_mem[1401] = 8'h00;
    red_mem[1402] = 8'h00;
    red_mem[1403] = 8'h00;
    red_mem[1404] = 8'h00;
    red_mem[1405] = 8'h00;
    red_mem[1406] = 8'h00;
    red_mem[1407] = 8'h00;
    red_mem[1408] = 8'h00;
    red_mem[1409] = 8'h00;
    red_mem[1410] = 8'h00;
    red_mem[1411] = 8'h00;
    red_mem[1412] = 8'h00;
    red_mem[1413] = 8'h00;
    red_mem[1414] = 8'h00;
    red_mem[1415] = 8'h00;
    red_mem[1416] = 8'h00;
    red_mem[1417] = 8'h00;
    red_mem[1418] = 8'h00;
    red_mem[1419] = 8'h00;
    red_mem[1420] = 8'h00;
    red_mem[1421] = 8'h00;
    red_mem[1422] = 8'h00;
    red_mem[1423] = 8'h00;
    red_mem[1424] = 8'h00;
    red_mem[1425] = 8'h00;
    red_mem[1426] = 8'h00;
    red_mem[1427] = 8'h00;
    red_mem[1428] = 8'h00;
    red_mem[1429] = 8'h00;
    red_mem[1430] = 8'h00;
    red_mem[1431] = 8'h00;
    red_mem[1432] = 8'h00;
    red_mem[1433] = 8'h00;
    red_mem[1434] = 8'h00;
    red_mem[1435] = 8'h00;
    red_mem[1436] = 8'h00;
    red_mem[1437] = 8'h00;
    red_mem[1438] = 8'h00;
    red_mem[1439] = 8'h00;
    red_mem[1440] = 8'h00;
    red_mem[1441] = 8'h00;
    red_mem[1442] = 8'h00;
    red_mem[1443] = 8'h00;
    red_mem[1444] = 8'h00;
    red_mem[1445] = 8'h00;
    red_mem[1446] = 8'h00;
    red_mem[1447] = 8'h00;
    red_mem[1448] = 8'h00;
    red_mem[1449] = 8'h00;
    red_mem[1450] = 8'h00;
    red_mem[1451] = 8'h00;
    red_mem[1452] = 8'h00;
    red_mem[1453] = 8'h00;
    red_mem[1454] = 8'h00;
    red_mem[1455] = 8'h00;
    red_mem[1456] = 8'h00;
    red_mem[1457] = 8'h00;
    red_mem[1458] = 8'h00;
    red_mem[1459] = 8'h00;
    red_mem[1460] = 8'h00;
    red_mem[1461] = 8'h00;
    red_mem[1462] = 8'h00;
    red_mem[1463] = 8'h00;
    red_mem[1464] = 8'h00;
    red_mem[1465] = 8'h00;
    red_mem[1466] = 8'h00;
    red_mem[1467] = 8'h00;
    red_mem[1468] = 8'h00;
    red_mem[1469] = 8'h00;
    red_mem[1470] = 8'h00;
    red_mem[1471] = 8'h00;
    red_mem[1472] = 8'h00;
    red_mem[1473] = 8'h00;
    red_mem[1474] = 8'h00;
    red_mem[1475] = 8'h00;
    red_mem[1476] = 8'h00;
    red_mem[1477] = 8'h00;
    red_mem[1478] = 8'h00;
    red_mem[1479] = 8'h00;
    red_mem[1480] = 8'h00;
    red_mem[1481] = 8'h00;
    red_mem[1482] = 8'h00;
    red_mem[1483] = 8'h00;
    red_mem[1484] = 8'h00;
    red_mem[1485] = 8'h00;
    red_mem[1486] = 8'h00;
    red_mem[1487] = 8'h00;
    red_mem[1488] = 8'h00;
    red_mem[1489] = 8'h00;
    red_mem[1490] = 8'h00;
    red_mem[1491] = 8'h00;
    red_mem[1492] = 8'h00;
    red_mem[1493] = 8'h00;
    red_mem[1494] = 8'h00;
    red_mem[1495] = 8'h00;
    red_mem[1496] = 8'h00;
    red_mem[1497] = 8'h00;
    red_mem[1498] = 8'h00;
    red_mem[1499] = 8'h00;
    red_mem[1500] = 8'h00;
    red_mem[1501] = 8'h00;
    red_mem[1502] = 8'h00;
    red_mem[1503] = 8'h00;
    red_mem[1504] = 8'h00;
    red_mem[1505] = 8'h00;
    red_mem[1506] = 8'h00;
    red_mem[1507] = 8'h00;
    red_mem[1508] = 8'h00;
    red_mem[1509] = 8'h00;
    red_mem[1510] = 8'h00;
    red_mem[1511] = 8'h00;
    red_mem[1512] = 8'h00;
    red_mem[1513] = 8'h00;
    red_mem[1514] = 8'h00;
    red_mem[1515] = 8'h00;
    red_mem[1516] = 8'h00;
    red_mem[1517] = 8'h00;
    red_mem[1518] = 8'h00;
    red_mem[1519] = 8'h00;
    red_mem[1520] = 8'h00;
    red_mem[1521] = 8'h00;
    red_mem[1522] = 8'h00;
    red_mem[1523] = 8'h00;
    red_mem[1524] = 8'h00;
    red_mem[1525] = 8'h00;
    red_mem[1526] = 8'h00;
    red_mem[1527] = 8'h00;
    red_mem[1528] = 8'h00;
    red_mem[1529] = 8'h00;
    red_mem[1530] = 8'h00;
    red_mem[1531] = 8'h00;
    red_mem[1532] = 8'h00;
    red_mem[1533] = 8'h00;
    red_mem[1534] = 8'h00;
    red_mem[1535] = 8'h00;
    red_mem[1536] = 8'h00;
    red_mem[1537] = 8'h00;
    red_mem[1538] = 8'h00;
    red_mem[1539] = 8'h00;
    red_mem[1540] = 8'h00;
    red_mem[1541] = 8'h00;
    red_mem[1542] = 8'h00;
    red_mem[1543] = 8'h00;
    red_mem[1544] = 8'h00;
    red_mem[1545] = 8'h00;
    red_mem[1546] = 8'h00;
    red_mem[1547] = 8'h00;
    red_mem[1548] = 8'h00;
    red_mem[1549] = 8'h00;
    red_mem[1550] = 8'h00;
    red_mem[1551] = 8'h00;
    red_mem[1552] = 8'h00;
    red_mem[1553] = 8'h00;
    red_mem[1554] = 8'h00;
    red_mem[1555] = 8'h00;
    red_mem[1556] = 8'h00;
    red_mem[1557] = 8'h00;
    red_mem[1558] = 8'h00;
    red_mem[1559] = 8'h00;
    red_mem[1560] = 8'h00;
    red_mem[1561] = 8'h00;
    red_mem[1562] = 8'h00;
    red_mem[1563] = 8'h00;
    red_mem[1564] = 8'h00;
    red_mem[1565] = 8'h00;
    red_mem[1566] = 8'h00;
    red_mem[1567] = 8'h00;
    red_mem[1568] = 8'h00;
    red_mem[1569] = 8'h00;
    red_mem[1570] = 8'h00;
    red_mem[1571] = 8'h00;
    red_mem[1572] = 8'h00;
    red_mem[1573] = 8'h00;
    red_mem[1574] = 8'h00;
    red_mem[1575] = 8'h00;
    red_mem[1576] = 8'h00;
    red_mem[1577] = 8'h00;
    red_mem[1578] = 8'h00;
    red_mem[1579] = 8'h00;
    red_mem[1580] = 8'h00;
    red_mem[1581] = 8'h00;
    red_mem[1582] = 8'h00;
    red_mem[1583] = 8'h00;
    red_mem[1584] = 8'h00;
    red_mem[1585] = 8'h00;
    red_mem[1586] = 8'h00;
    red_mem[1587] = 8'h00;
    red_mem[1588] = 8'h00;
    red_mem[1589] = 8'h00;
    red_mem[1590] = 8'h00;
    red_mem[1591] = 8'h00;
    red_mem[1592] = 8'h00;
    red_mem[1593] = 8'h00;
    red_mem[1594] = 8'h00;
    red_mem[1595] = 8'h00;
    red_mem[1596] = 8'h00;
    red_mem[1597] = 8'h00;
    red_mem[1598] = 8'h00;
    red_mem[1599] = 8'h00;
    red_mem[1600] = 8'h00;
    red_mem[1601] = 8'h00;
    red_mem[1602] = 8'h00;
    red_mem[1603] = 8'h00;
    red_mem[1604] = 8'h00;
    red_mem[1605] = 8'h00;
    red_mem[1606] = 8'h00;
    red_mem[1607] = 8'h00;
    red_mem[1608] = 8'h00;
    red_mem[1609] = 8'h00;
    red_mem[1610] = 8'h00;
    red_mem[1611] = 8'h00;
    red_mem[1612] = 8'h00;
    red_mem[1613] = 8'h00;
    red_mem[1614] = 8'h00;
    red_mem[1615] = 8'h00;
    red_mem[1616] = 8'h00;
    red_mem[1617] = 8'h00;
    red_mem[1618] = 8'h00;
    red_mem[1619] = 8'h00;
    red_mem[1620] = 8'h00;
    red_mem[1621] = 8'h00;
    red_mem[1622] = 8'h00;
    red_mem[1623] = 8'h00;
    red_mem[1624] = 8'h00;
    red_mem[1625] = 8'h00;
    red_mem[1626] = 8'h00;
    red_mem[1627] = 8'h00;
    red_mem[1628] = 8'h00;
    red_mem[1629] = 8'h00;
    red_mem[1630] = 8'h00;
    red_mem[1631] = 8'h00;
    red_mem[1632] = 8'h00;
    red_mem[1633] = 8'h00;
    red_mem[1634] = 8'h00;
    red_mem[1635] = 8'h00;
    red_mem[1636] = 8'h00;
    red_mem[1637] = 8'h00;
    red_mem[1638] = 8'h00;
    red_mem[1639] = 8'h00;
    red_mem[1640] = 8'h00;
    red_mem[1641] = 8'h00;
    red_mem[1642] = 8'h00;
    red_mem[1643] = 8'h00;
    red_mem[1644] = 8'h00;
    red_mem[1645] = 8'h00;
    red_mem[1646] = 8'h00;
    red_mem[1647] = 8'h00;
    red_mem[1648] = 8'h00;
    red_mem[1649] = 8'h00;
    red_mem[1650] = 8'h00;
    red_mem[1651] = 8'h00;
    red_mem[1652] = 8'h00;
    red_mem[1653] = 8'h00;
    red_mem[1654] = 8'h00;
    red_mem[1655] = 8'h00;
    red_mem[1656] = 8'h00;
    red_mem[1657] = 8'h00;
    red_mem[1658] = 8'h00;
    red_mem[1659] = 8'h00;
    red_mem[1660] = 8'h00;
    red_mem[1661] = 8'h00;
    red_mem[1662] = 8'h00;
    red_mem[1663] = 8'h00;
    red_mem[1664] = 8'h00;
    red_mem[1665] = 8'h00;
    red_mem[1666] = 8'h00;
    red_mem[1667] = 8'h00;
    red_mem[1668] = 8'h00;
    red_mem[1669] = 8'h00;
    red_mem[1670] = 8'h00;
    red_mem[1671] = 8'h00;
    red_mem[1672] = 8'h00;
    red_mem[1673] = 8'h00;
    red_mem[1674] = 8'h00;
    red_mem[1675] = 8'h00;
    red_mem[1676] = 8'h00;
    red_mem[1677] = 8'h00;
    red_mem[1678] = 8'h00;
    red_mem[1679] = 8'h00;
    red_mem[1680] = 8'h00;
    red_mem[1681] = 8'h00;
    red_mem[1682] = 8'h00;
    red_mem[1683] = 8'h00;
    red_mem[1684] = 8'h00;
    red_mem[1685] = 8'h00;
    red_mem[1686] = 8'h00;
    red_mem[1687] = 8'h00;
    red_mem[1688] = 8'h00;
    red_mem[1689] = 8'h00;
    red_mem[1690] = 8'h00;
    red_mem[1691] = 8'h00;
    red_mem[1692] = 8'h00;
    red_mem[1693] = 8'h00;
    red_mem[1694] = 8'h00;
    red_mem[1695] = 8'h00;
    red_mem[1696] = 8'h00;
    red_mem[1697] = 8'h00;
    red_mem[1698] = 8'h00;
    red_mem[1699] = 8'h00;
    red_mem[1700] = 8'h00;
    red_mem[1701] = 8'h00;
    red_mem[1702] = 8'h00;
    red_mem[1703] = 8'h00;
    red_mem[1704] = 8'h00;
    red_mem[1705] = 8'h00;
    red_mem[1706] = 8'h00;
    red_mem[1707] = 8'h00;
    red_mem[1708] = 8'h00;
    red_mem[1709] = 8'h00;
    red_mem[1710] = 8'h00;
    red_mem[1711] = 8'h00;
    red_mem[1712] = 8'h00;
    red_mem[1713] = 8'h00;
    red_mem[1714] = 8'h00;
    red_mem[1715] = 8'h00;
    red_mem[1716] = 8'h00;
    red_mem[1717] = 8'h00;
    red_mem[1718] = 8'h00;
    red_mem[1719] = 8'h00;
    red_mem[1720] = 8'h00;
    red_mem[1721] = 8'h00;
    red_mem[1722] = 8'h00;
    red_mem[1723] = 8'h00;
    red_mem[1724] = 8'h00;
    red_mem[1725] = 8'h00;
    red_mem[1726] = 8'h00;
    red_mem[1727] = 8'h00;
    red_mem[1728] = 8'h00;
    red_mem[1729] = 8'h00;
    red_mem[1730] = 8'h00;
    red_mem[1731] = 8'h00;
    red_mem[1732] = 8'h00;
    red_mem[1733] = 8'h00;
    red_mem[1734] = 8'h00;
    red_mem[1735] = 8'h00;
    red_mem[1736] = 8'h00;
    red_mem[1737] = 8'h00;
    red_mem[1738] = 8'h00;
    red_mem[1739] = 8'h00;
    red_mem[1740] = 8'h00;
    red_mem[1741] = 8'h00;
    red_mem[1742] = 8'h00;
    red_mem[1743] = 8'h00;
    red_mem[1744] = 8'h00;
    red_mem[1745] = 8'h00;
    red_mem[1746] = 8'h00;
    red_mem[1747] = 8'h00;
    red_mem[1748] = 8'h00;
    red_mem[1749] = 8'h00;
    red_mem[1750] = 8'h00;
    red_mem[1751] = 8'h00;
    red_mem[1752] = 8'h00;
    red_mem[1753] = 8'h00;
    red_mem[1754] = 8'h00;
    red_mem[1755] = 8'h00;
    red_mem[1756] = 8'h00;
    red_mem[1757] = 8'h00;
    red_mem[1758] = 8'h00;
    red_mem[1759] = 8'h00;
    red_mem[1760] = 8'h00;
    red_mem[1761] = 8'h00;
    red_mem[1762] = 8'h00;
    red_mem[1763] = 8'h00;
    red_mem[1764] = 8'h00;
    red_mem[1765] = 8'h00;
    red_mem[1766] = 8'h00;
    red_mem[1767] = 8'h00;
    red_mem[1768] = 8'h00;
    red_mem[1769] = 8'h00;
    red_mem[1770] = 8'h00;
    red_mem[1771] = 8'h00;
    red_mem[1772] = 8'h00;
    red_mem[1773] = 8'h00;
    red_mem[1774] = 8'h00;
    red_mem[1775] = 8'h00;
    red_mem[1776] = 8'h00;
    red_mem[1777] = 8'h00;
    red_mem[1778] = 8'h00;
    red_mem[1779] = 8'h00;
    red_mem[1780] = 8'h00;
    red_mem[1781] = 8'h00;
    red_mem[1782] = 8'h00;
    red_mem[1783] = 8'h00;
    red_mem[1784] = 8'h00;
    red_mem[1785] = 8'h00;
    red_mem[1786] = 8'h00;
    red_mem[1787] = 8'h00;
    red_mem[1788] = 8'h00;
    red_mem[1789] = 8'h00;
    red_mem[1790] = 8'h00;
    red_mem[1791] = 8'h00;
    red_mem[1792] = 8'h00;
    red_mem[1793] = 8'h00;
    red_mem[1794] = 8'h00;
    red_mem[1795] = 8'h00;
    red_mem[1796] = 8'h00;
    red_mem[1797] = 8'h00;
    red_mem[1798] = 8'h00;
    red_mem[1799] = 8'h00;
    red_mem[1800] = 8'h00;
    red_mem[1801] = 8'h00;
    red_mem[1802] = 8'h00;
    red_mem[1803] = 8'h00;
    red_mem[1804] = 8'h00;
    red_mem[1805] = 8'h00;
    red_mem[1806] = 8'h00;
    red_mem[1807] = 8'h00;
    red_mem[1808] = 8'h00;
    red_mem[1809] = 8'h00;
    red_mem[1810] = 8'h00;
    red_mem[1811] = 8'h00;
    red_mem[1812] = 8'h00;
    red_mem[1813] = 8'h00;
    red_mem[1814] = 8'h00;
    red_mem[1815] = 8'h00;
    red_mem[1816] = 8'h00;
    red_mem[1817] = 8'h00;
    red_mem[1818] = 8'h00;
    red_mem[1819] = 8'h00;
    red_mem[1820] = 8'h00;
    red_mem[1821] = 8'h00;
    red_mem[1822] = 8'h00;
    red_mem[1823] = 8'h00;
    red_mem[1824] = 8'h00;
    red_mem[1825] = 8'h00;
    red_mem[1826] = 8'h00;
    red_mem[1827] = 8'h00;
    red_mem[1828] = 8'h00;
    red_mem[1829] = 8'h00;
    red_mem[1830] = 8'h00;
    red_mem[1831] = 8'h00;
    red_mem[1832] = 8'h00;
    red_mem[1833] = 8'h00;
    red_mem[1834] = 8'h00;
    red_mem[1835] = 8'h00;
    red_mem[1836] = 8'h00;
    red_mem[1837] = 8'h00;
    red_mem[1838] = 8'h00;
    red_mem[1839] = 8'h00;
    red_mem[1840] = 8'h00;
    red_mem[1841] = 8'h00;
    red_mem[1842] = 8'h00;
    red_mem[1843] = 8'h00;
    red_mem[1844] = 8'h00;
    red_mem[1845] = 8'h00;
    red_mem[1846] = 8'h00;
    red_mem[1847] = 8'h00;
    red_mem[1848] = 8'h00;
    red_mem[1849] = 8'h00;
    red_mem[1850] = 8'h00;
    red_mem[1851] = 8'h00;
    red_mem[1852] = 8'h00;
    red_mem[1853] = 8'h00;
    red_mem[1854] = 8'h00;
    red_mem[1855] = 8'h00;
    red_mem[1856] = 8'h00;
    red_mem[1857] = 8'h00;
    red_mem[1858] = 8'h00;
    red_mem[1859] = 8'h00;
    red_mem[1860] = 8'h00;
    red_mem[1861] = 8'h00;
    red_mem[1862] = 8'h00;
    red_mem[1863] = 8'h00;
    red_mem[1864] = 8'h00;
    red_mem[1865] = 8'h00;
    red_mem[1866] = 8'h00;
    red_mem[1867] = 8'h00;
    red_mem[1868] = 8'h00;
    red_mem[1869] = 8'h00;
    red_mem[1870] = 8'h00;
    red_mem[1871] = 8'h00;
    red_mem[1872] = 8'h00;
    red_mem[1873] = 8'h00;
    red_mem[1874] = 8'h00;
    red_mem[1875] = 8'h00;
    red_mem[1876] = 8'h00;
    red_mem[1877] = 8'h00;
    red_mem[1878] = 8'h00;
    red_mem[1879] = 8'h00;
    red_mem[1880] = 8'h00;
    red_mem[1881] = 8'h00;
    red_mem[1882] = 8'h00;
    red_mem[1883] = 8'h00;
    red_mem[1884] = 8'h00;
    red_mem[1885] = 8'h00;
    red_mem[1886] = 8'h00;
    red_mem[1887] = 8'h00;
    red_mem[1888] = 8'h00;
    red_mem[1889] = 8'h00;
    red_mem[1890] = 8'h00;
    red_mem[1891] = 8'h00;
    red_mem[1892] = 8'h00;
    red_mem[1893] = 8'h00;
    red_mem[1894] = 8'h00;
    red_mem[1895] = 8'h00;
    red_mem[1896] = 8'h00;
    red_mem[1897] = 8'h00;
    red_mem[1898] = 8'h00;
    red_mem[1899] = 8'h00;
    red_mem[1900] = 8'h00;
    red_mem[1901] = 8'h00;
    red_mem[1902] = 8'h00;
    red_mem[1903] = 8'h00;
    red_mem[1904] = 8'h00;
    red_mem[1905] = 8'h00;
    red_mem[1906] = 8'h00;
    red_mem[1907] = 8'h00;
    red_mem[1908] = 8'h00;
    red_mem[1909] = 8'h00;
    red_mem[1910] = 8'h00;
    red_mem[1911] = 8'h00;
    red_mem[1912] = 8'h00;
    red_mem[1913] = 8'h00;
    red_mem[1914] = 8'h00;
    red_mem[1915] = 8'h00;
    red_mem[1916] = 8'h00;
    red_mem[1917] = 8'h00;
    red_mem[1918] = 8'h00;
    red_mem[1919] = 8'h00;
    red_mem[1920] = 8'h00;
    red_mem[1921] = 8'h00;
    red_mem[1922] = 8'h00;
    red_mem[1923] = 8'h00;
    red_mem[1924] = 8'h00;
    red_mem[1925] = 8'h00;
    red_mem[1926] = 8'h00;
    red_mem[1927] = 8'h00;
    red_mem[1928] = 8'h00;
    red_mem[1929] = 8'h00;
    red_mem[1930] = 8'h00;
    red_mem[1931] = 8'h00;
    red_mem[1932] = 8'h00;
    red_mem[1933] = 8'h00;
    red_mem[1934] = 8'h00;
    red_mem[1935] = 8'h00;
    red_mem[1936] = 8'h00;
    red_mem[1937] = 8'h00;
    red_mem[1938] = 8'h00;
    red_mem[1939] = 8'h00;
    red_mem[1940] = 8'h00;
    red_mem[1941] = 8'h00;
    red_mem[1942] = 8'h00;
    red_mem[1943] = 8'h00;
    red_mem[1944] = 8'h00;
    red_mem[1945] = 8'h00;
    red_mem[1946] = 8'h00;
    red_mem[1947] = 8'h00;
    red_mem[1948] = 8'h00;
    red_mem[1949] = 8'h00;
    red_mem[1950] = 8'h00;
    red_mem[1951] = 8'h00;
    red_mem[1952] = 8'h00;
    red_mem[1953] = 8'h00;
    red_mem[1954] = 8'h00;
    red_mem[1955] = 8'h00;
    red_mem[1956] = 8'h00;
    red_mem[1957] = 8'h00;
    red_mem[1958] = 8'h00;
    red_mem[1959] = 8'h00;
    red_mem[1960] = 8'h00;
    red_mem[1961] = 8'h00;
    red_mem[1962] = 8'h00;
    red_mem[1963] = 8'h00;
    red_mem[1964] = 8'h00;
    red_mem[1965] = 8'h00;
    red_mem[1966] = 8'h00;
    red_mem[1967] = 8'h00;
    red_mem[1968] = 8'h00;
    red_mem[1969] = 8'h00;
    red_mem[1970] = 8'h00;
    red_mem[1971] = 8'h00;
    red_mem[1972] = 8'h00;
    red_mem[1973] = 8'h00;
    red_mem[1974] = 8'h00;
    red_mem[1975] = 8'h00;
    red_mem[1976] = 8'h00;
    red_mem[1977] = 8'h00;
    red_mem[1978] = 8'h00;
    red_mem[1979] = 8'h00;
    red_mem[1980] = 8'h00;
    red_mem[1981] = 8'h00;
    red_mem[1982] = 8'h00;
    red_mem[1983] = 8'h00;
    red_mem[1984] = 8'h00;
    red_mem[1985] = 8'h00;
    red_mem[1986] = 8'h00;
    red_mem[1987] = 8'h00;
    red_mem[1988] = 8'h00;
    red_mem[1989] = 8'h00;
    red_mem[1990] = 8'h00;
    red_mem[1991] = 8'h00;
    red_mem[1992] = 8'h00;
    red_mem[1993] = 8'h00;
    red_mem[1994] = 8'h00;
    red_mem[1995] = 8'h00;
    red_mem[1996] = 8'h00;
    red_mem[1997] = 8'h00;
    red_mem[1998] = 8'h00;
    red_mem[1999] = 8'h00;
    red_mem[2000] = 8'h00;
    red_mem[2001] = 8'h00;
    red_mem[2002] = 8'h00;
    red_mem[2003] = 8'h00;
    red_mem[2004] = 8'h00;
    red_mem[2005] = 8'h00;
    red_mem[2006] = 8'h00;
    red_mem[2007] = 8'h00;
    red_mem[2008] = 8'h00;
    red_mem[2009] = 8'h00;
    red_mem[2010] = 8'h00;
    red_mem[2011] = 8'h00;
    red_mem[2012] = 8'h00;
    red_mem[2013] = 8'h00;
    red_mem[2014] = 8'h00;
    red_mem[2015] = 8'h00;
    red_mem[2016] = 8'h00;
    red_mem[2017] = 8'h00;
    red_mem[2018] = 8'h00;
    red_mem[2019] = 8'h00;
    red_mem[2020] = 8'h00;
    red_mem[2021] = 8'h00;
    red_mem[2022] = 8'h00;
    red_mem[2023] = 8'h00;
    red_mem[2024] = 8'h00;
    red_mem[2025] = 8'h00;
    red_mem[2026] = 8'h00;
    red_mem[2027] = 8'h00;
    red_mem[2028] = 8'h00;
    red_mem[2029] = 8'h00;
    red_mem[2030] = 8'h00;
    red_mem[2031] = 8'h00;
    red_mem[2032] = 8'h00;
    red_mem[2033] = 8'h00;
    red_mem[2034] = 8'h00;
    red_mem[2035] = 8'h00;
    red_mem[2036] = 8'h00;
    red_mem[2037] = 8'h00;
    red_mem[2038] = 8'h00;
    red_mem[2039] = 8'h00;
    red_mem[2040] = 8'h00;
    red_mem[2041] = 8'h00;
    red_mem[2042] = 8'h00;
    red_mem[2043] = 8'h00;
    red_mem[2044] = 8'h00;
    red_mem[2045] = 8'h00;
    red_mem[2046] = 8'h00;
    red_mem[2047] = 8'h00;
    green_mem[0] = 8'h00;
    green_mem[1] = 8'h00;
    green_mem[2] = 8'h00;
    green_mem[3] = 8'h00;
    green_mem[4] = 8'h00;
    green_mem[5] = 8'h00;
    green_mem[6] = 8'h00;
    green_mem[7] = 8'h00;
    green_mem[8] = 8'h00;
    green_mem[9] = 8'h00;
    green_mem[10] = 8'h00;
    green_mem[11] = 8'h00;
    green_mem[12] = 8'h00;
    green_mem[13] = 8'h00;
    green_mem[14] = 8'h00;
    green_mem[15] = 8'h00;
    green_mem[16] = 8'h00;
    green_mem[17] = 8'h00;
    green_mem[18] = 8'h00;
    green_mem[19] = 8'h00;
    green_mem[20] = 8'h00;
    green_mem[21] = 8'h00;
    green_mem[22] = 8'h00;
    green_mem[23] = 8'h00;
    green_mem[24] = 8'h00;
    green_mem[25] = 8'h00;
    green_mem[26] = 8'h00;
    green_mem[27] = 8'h00;
    green_mem[28] = 8'h00;
    green_mem[29] = 8'h00;
    green_mem[30] = 8'h00;
    green_mem[31] = 8'h00;
    green_mem[32] = 8'h00;
    green_mem[33] = 8'h00;
    green_mem[34] = 8'h00;
    green_mem[35] = 8'h00;
    green_mem[36] = 8'h00;
    green_mem[37] = 8'h00;
    green_mem[38] = 8'h00;
    green_mem[39] = 8'h00;
    green_mem[40] = 8'h00;
    green_mem[41] = 8'h00;
    green_mem[42] = 8'h00;
    green_mem[43] = 8'h00;
    green_mem[44] = 8'h00;
    green_mem[45] = 8'h00;
    green_mem[46] = 8'h00;
    green_mem[47] = 8'h00;
    green_mem[48] = 8'h00;
    green_mem[49] = 8'h00;
    green_mem[50] = 8'h00;
    green_mem[51] = 8'h00;
    green_mem[52] = 8'h00;
    green_mem[53] = 8'h00;
    green_mem[54] = 8'h00;
    green_mem[55] = 8'h00;
    green_mem[56] = 8'h00;
    green_mem[57] = 8'h00;
    green_mem[58] = 8'h00;
    green_mem[59] = 8'h00;
    green_mem[60] = 8'h00;
    green_mem[61] = 8'h00;
    green_mem[62] = 8'h00;
    green_mem[63] = 8'h00;
    green_mem[64] = 8'h00;
    green_mem[65] = 8'h00;
    green_mem[66] = 8'h00;
    green_mem[67] = 8'h00;
    green_mem[68] = 8'h00;
    green_mem[69] = 8'h00;
    green_mem[70] = 8'h00;
    green_mem[71] = 8'h00;
    green_mem[72] = 8'h00;
    green_mem[73] = 8'h00;
    green_mem[74] = 8'h00;
    green_mem[75] = 8'h00;
    green_mem[76] = 8'h00;
    green_mem[77] = 8'h00;
    green_mem[78] = 8'h00;
    green_mem[79] = 8'h00;
    green_mem[80] = 8'h00;
    green_mem[81] = 8'h00;
    green_mem[82] = 8'h00;
    green_mem[83] = 8'h00;
    green_mem[84] = 8'h00;
    green_mem[85] = 8'h00;
    green_mem[86] = 8'h00;
    green_mem[87] = 8'h00;
    green_mem[88] = 8'h00;
    green_mem[89] = 8'h00;
    green_mem[90] = 8'h00;
    green_mem[91] = 8'h00;
    green_mem[92] = 8'h00;
    green_mem[93] = 8'h00;
    green_mem[94] = 8'h00;
    green_mem[95] = 8'h00;
    green_mem[96] = 8'h00;
    green_mem[97] = 8'h00;
    green_mem[98] = 8'h00;
    green_mem[99] = 8'h00;
    green_mem[100] = 8'h00;
    green_mem[101] = 8'h00;
    green_mem[102] = 8'h00;
    green_mem[103] = 8'h00;
    green_mem[104] = 8'h00;
    green_mem[105] = 8'h00;
    green_mem[106] = 8'h00;
    green_mem[107] = 8'h00;
    green_mem[108] = 8'h00;
    green_mem[109] = 8'h00;
    green_mem[110] = 8'h00;
    green_mem[111] = 8'h00;
    green_mem[112] = 8'h00;
    green_mem[113] = 8'h00;
    green_mem[114] = 8'h00;
    green_mem[115] = 8'h00;
    green_mem[116] = 8'h00;
    green_mem[117] = 8'h00;
    green_mem[118] = 8'h00;
    green_mem[119] = 8'h00;
    green_mem[120] = 8'h00;
    green_mem[121] = 8'h00;
    green_mem[122] = 8'h00;
    green_mem[123] = 8'h00;
    green_mem[124] = 8'h00;
    green_mem[125] = 8'h00;
    green_mem[126] = 8'h00;
    green_mem[127] = 8'h00;
    green_mem[128] = 8'h00;
    green_mem[129] = 8'h00;
    green_mem[130] = 8'h00;
    green_mem[131] = 8'h00;
    green_mem[132] = 8'h00;
    green_mem[133] = 8'h00;
    green_mem[134] = 8'h00;
    green_mem[135] = 8'h00;
    green_mem[136] = 8'h00;
    green_mem[137] = 8'h00;
    green_mem[138] = 8'h00;
    green_mem[139] = 8'h00;
    green_mem[140] = 8'h00;
    green_mem[141] = 8'h00;
    green_mem[142] = 8'h00;
    green_mem[143] = 8'h00;
    green_mem[144] = 8'h00;
    green_mem[145] = 8'h00;
    green_mem[146] = 8'h00;
    green_mem[147] = 8'h00;
    green_mem[148] = 8'h00;
    green_mem[149] = 8'h00;
    green_mem[150] = 8'h00;
    green_mem[151] = 8'h00;
    green_mem[152] = 8'h00;
    green_mem[153] = 8'h00;
    green_mem[154] = 8'h00;
    green_mem[155] = 8'h00;
    green_mem[156] = 8'h00;
    green_mem[157] = 8'h00;
    green_mem[158] = 8'h00;
    green_mem[159] = 8'h00;
    green_mem[160] = 8'h00;
    green_mem[161] = 8'h00;
    green_mem[162] = 8'h00;
    green_mem[163] = 8'h00;
    green_mem[164] = 8'h00;
    green_mem[165] = 8'h00;
    green_mem[166] = 8'h00;
    green_mem[167] = 8'h00;
    green_mem[168] = 8'h00;
    green_mem[169] = 8'h00;
    green_mem[170] = 8'h00;
    green_mem[171] = 8'h00;
    green_mem[172] = 8'h00;
    green_mem[173] = 8'h00;
    green_mem[174] = 8'h00;
    green_mem[175] = 8'h00;
    green_mem[176] = 8'h00;
    green_mem[177] = 8'h00;
    green_mem[178] = 8'h00;
    green_mem[179] = 8'h00;
    green_mem[180] = 8'h00;
    green_mem[181] = 8'h00;
    green_mem[182] = 8'h00;
    green_mem[183] = 8'h00;
    green_mem[184] = 8'h00;
    green_mem[185] = 8'h00;
    green_mem[186] = 8'h00;
    green_mem[187] = 8'h00;
    green_mem[188] = 8'h00;
    green_mem[189] = 8'h00;
    green_mem[190] = 8'h00;
    green_mem[191] = 8'h00;
    green_mem[192] = 8'h00;
    green_mem[193] = 8'h00;
    green_mem[194] = 8'h00;
    green_mem[195] = 8'h00;
    green_mem[196] = 8'h00;
    green_mem[197] = 8'h00;
    green_mem[198] = 8'h00;
    green_mem[199] = 8'h00;
    green_mem[200] = 8'h00;
    green_mem[201] = 8'h00;
    green_mem[202] = 8'h00;
    green_mem[203] = 8'h00;
    green_mem[204] = 8'h00;
    green_mem[205] = 8'h00;
    green_mem[206] = 8'h00;
    green_mem[207] = 8'h00;
    green_mem[208] = 8'h00;
    green_mem[209] = 8'h00;
    green_mem[210] = 8'h00;
    green_mem[211] = 8'h00;
    green_mem[212] = 8'h00;
    green_mem[213] = 8'h00;
    green_mem[214] = 8'h00;
    green_mem[215] = 8'h00;
    green_mem[216] = 8'h00;
    green_mem[217] = 8'h00;
    green_mem[218] = 8'h00;
    green_mem[219] = 8'h00;
    green_mem[220] = 8'h00;
    green_mem[221] = 8'h00;
    green_mem[222] = 8'h00;
    green_mem[223] = 8'h00;
    green_mem[224] = 8'h00;
    green_mem[225] = 8'h00;
    green_mem[226] = 8'h00;
    green_mem[227] = 8'h00;
    green_mem[228] = 8'h00;
    green_mem[229] = 8'h00;
    green_mem[230] = 8'h00;
    green_mem[231] = 8'h00;
    green_mem[232] = 8'h00;
    green_mem[233] = 8'h00;
    green_mem[234] = 8'h00;
    green_mem[235] = 8'h00;
    green_mem[236] = 8'h00;
    green_mem[237] = 8'h00;
    green_mem[238] = 8'h00;
    green_mem[239] = 8'h00;
    green_mem[240] = 8'h00;
    green_mem[241] = 8'h00;
    green_mem[242] = 8'h00;
    green_mem[243] = 8'h00;
    green_mem[244] = 8'h00;
    green_mem[245] = 8'h00;
    green_mem[246] = 8'h00;
    green_mem[247] = 8'h00;
    green_mem[248] = 8'h00;
    green_mem[249] = 8'h00;
    green_mem[250] = 8'h00;
    green_mem[251] = 8'h00;
    green_mem[252] = 8'h00;
    green_mem[253] = 8'h00;
    green_mem[254] = 8'h00;
    green_mem[255] = 8'h00;
    green_mem[256] = 8'h00;
    green_mem[257] = 8'h00;
    green_mem[258] = 8'h00;
    green_mem[259] = 8'h00;
    green_mem[260] = 8'h00;
    green_mem[261] = 8'h00;
    green_mem[262] = 8'h00;
    green_mem[263] = 8'h00;
    green_mem[264] = 8'h10;
    green_mem[265] = 8'h00;
    green_mem[266] = 8'h00;
    green_mem[267] = 8'h00;
    green_mem[268] = 8'h00;
    green_mem[269] = 8'h00;
    green_mem[270] = 8'h00;
    green_mem[271] = 8'h00;
    green_mem[272] = 8'h00;
    green_mem[273] = 8'h00;
    green_mem[274] = 8'h00;
    green_mem[275] = 8'h00;
    green_mem[276] = 8'h00;
    green_mem[277] = 8'h00;
    green_mem[278] = 8'h00;
    green_mem[279] = 8'hd8;
    green_mem[280] = 8'hfd;
    green_mem[281] = 8'h03;
    green_mem[282] = 8'h00;
    green_mem[283] = 8'h00;
    green_mem[284] = 8'h00;
    green_mem[285] = 8'h00;
    green_mem[286] = 8'h00;
    green_mem[287] = 8'h00;
    green_mem[288] = 8'h00;
    green_mem[289] = 8'h00;
    green_mem[290] = 8'h00;
    green_mem[291] = 8'h00;
    green_mem[292] = 8'h00;
    green_mem[293] = 8'h00;
    green_mem[294] = 8'hb8;
    green_mem[295] = 8'hff;
    green_mem[296] = 8'hff;
    green_mem[297] = 8'h3b;
    green_mem[298] = 8'h00;
    green_mem[299] = 8'h00;
    green_mem[300] = 8'h00;
    green_mem[301] = 8'h00;
    green_mem[302] = 8'h00;
    green_mem[303] = 8'h00;
    green_mem[304] = 8'h00;
    green_mem[305] = 8'h00;
    green_mem[306] = 8'h00;
    green_mem[307] = 8'h00;
    green_mem[308] = 8'h00;
    green_mem[309] = 8'h00;
    green_mem[310] = 8'hfc;
    green_mem[311] = 8'hff;
    green_mem[312] = 8'hff;
    green_mem[313] = 8'hfb;
    green_mem[314] = 8'h03;
    green_mem[315] = 8'h00;
    green_mem[316] = 8'h00;
    green_mem[317] = 8'h00;
    green_mem[318] = 8'h00;
    green_mem[319] = 8'h00;
    green_mem[320] = 8'h00;
    green_mem[321] = 8'h00;
    green_mem[322] = 8'h00;
    green_mem[323] = 8'h00;
    green_mem[324] = 8'h00;
    green_mem[325] = 8'hc0;
    green_mem[326] = 8'hff;
    green_mem[327] = 8'hff;
    green_mem[328] = 8'hff;
    green_mem[329] = 8'hff;
    green_mem[330] = 8'h03;
    green_mem[331] = 8'h00;
    green_mem[332] = 8'h00;
    green_mem[333] = 8'h00;
    green_mem[334] = 8'h00;
    green_mem[335] = 8'h00;
    green_mem[336] = 8'h00;
    green_mem[337] = 8'h00;
    green_mem[338] = 8'h00;
    green_mem[339] = 8'h00;
    green_mem[340] = 8'h00;
    green_mem[341] = 8'he0;
    green_mem[342] = 8'hff;
    green_mem[343] = 8'hff;
    green_mem[344] = 8'hff;
    green_mem[345] = 8'hff;
    green_mem[346] = 8'h17;
    green_mem[347] = 8'h00;
    green_mem[348] = 8'h00;
    green_mem[349] = 8'h00;
    green_mem[350] = 8'h00;
    green_mem[351] = 8'h00;
    green_mem[352] = 8'h00;
    green_mem[353] = 8'h00;
    green_mem[354] = 8'h00;
    green_mem[355] = 8'h00;
    green_mem[356] = 8'h00;
    green_mem[357] = 8'hfc;
    green_mem[358] = 8'hff;
    green_mem[359] = 8'hff;
    green_mem[360] = 8'hff;
    green_mem[361] = 8'hff;
    green_mem[362] = 8'h3f;
    green_mem[363] = 8'h00;
    green_mem[364] = 8'h00;
    green_mem[365] = 8'h00;
    green_mem[366] = 8'h00;
    green_mem[367] = 8'h00;
    green_mem[368] = 8'h00;
    green_mem[369] = 8'h00;
    green_mem[370] = 8'h00;
    green_mem[371] = 8'h00;
    green_mem[372] = 8'h00;
    green_mem[373] = 8'hfc;
    green_mem[374] = 8'hff;
    green_mem[375] = 8'hff;
    green_mem[376] = 8'hff;
    green_mem[377] = 8'hff;
    green_mem[378] = 8'h3f;
    green_mem[379] = 8'h00;
    green_mem[380] = 8'h00;
    green_mem[381] = 8'h00;
    green_mem[382] = 8'h00;
    green_mem[383] = 8'h00;
    green_mem[384] = 8'h00;
    green_mem[385] = 8'h00;
    green_mem[386] = 8'h00;
    green_mem[387] = 8'h00;
    green_mem[388] = 8'hc0;
    green_mem[389] = 8'hff;
    green_mem[390] = 8'hff;
    green_mem[391] = 8'hff;
    green_mem[392] = 8'hff;
    green_mem[393] = 8'hff;
    green_mem[394] = 8'hff;
    green_mem[395] = 8'h07;
    green_mem[396] = 8'h00;
    green_mem[397] = 8'h00;
    green_mem[398] = 8'h00;
    green_mem[399] = 8'h00;
    green_mem[400] = 8'h00;
    green_mem[401] = 8'h00;
    green_mem[402] = 8'h00;
    green_mem[403] = 8'h00;
    green_mem[404] = 8'hc0;
    green_mem[405] = 8'hff;
    green_mem[406] = 8'hff;
    green_mem[407] = 8'hff;
    green_mem[408] = 8'hff;
    green_mem[409] = 8'hff;
    green_mem[410] = 8'hff;
    green_mem[411] = 8'h0f;
    green_mem[412] = 8'h00;
    green_mem[413] = 8'h00;
    green_mem[414] = 8'h00;
    green_mem[415] = 8'h00;
    green_mem[416] = 8'h00;
    green_mem[417] = 8'h00;
    green_mem[418] = 8'h00;
    green_mem[419] = 8'h00;
    green_mem[420] = 8'hf8;
    green_mem[421] = 8'hff;
    green_mem[422] = 8'hff;
    green_mem[423] = 8'hff;
    green_mem[424] = 8'hff;
    green_mem[425] = 8'hff;
    green_mem[426] = 8'hff;
    green_mem[427] = 8'h0f;
    green_mem[428] = 8'h00;
    green_mem[429] = 8'h00;
    green_mem[430] = 8'h00;
    green_mem[431] = 8'h00;
    green_mem[432] = 8'h00;
    green_mem[433] = 8'h00;
    green_mem[434] = 8'h00;
    green_mem[435] = 8'h00;
    green_mem[436] = 8'hf8;
    green_mem[437] = 8'hff;
    green_mem[438] = 8'hbf;
    green_mem[439] = 8'hff;
    green_mem[440] = 8'hff;
    green_mem[441] = 8'hff;
    green_mem[442] = 8'hff;
    green_mem[443] = 8'h3f;
    green_mem[444] = 8'h00;
    green_mem[445] = 8'h00;
    green_mem[446] = 8'h00;
    green_mem[447] = 8'h00;
    green_mem[448] = 8'h00;
    green_mem[449] = 8'h00;
    green_mem[450] = 8'h00;
    green_mem[451] = 8'h00;
    green_mem[452] = 8'hf8;
    green_mem[453] = 8'hff;
    green_mem[454] = 8'hff;
    green_mem[455] = 8'hff;
    green_mem[456] = 8'hff;
    green_mem[457] = 8'hff;
    green_mem[458] = 8'hff;
    green_mem[459] = 8'h7f;
    green_mem[460] = 8'h00;
    green_mem[461] = 8'h00;
    green_mem[462] = 8'h00;
    green_mem[463] = 8'h00;
    green_mem[464] = 8'h00;
    green_mem[465] = 8'h00;
    green_mem[466] = 8'h00;
    green_mem[467] = 8'h00;
    green_mem[468] = 8'hfe;
    green_mem[469] = 8'hff;
    green_mem[470] = 8'hff;
    green_mem[471] = 8'hff;
    green_mem[472] = 8'hff;
    green_mem[473] = 8'hff;
    green_mem[474] = 8'hff;
    green_mem[475] = 8'hff;
    green_mem[476] = 8'h01;
    green_mem[477] = 8'h00;
    green_mem[478] = 8'h00;
    green_mem[479] = 8'h00;
    green_mem[480] = 8'h00;
    green_mem[481] = 8'h00;
    green_mem[482] = 8'h00;
    green_mem[483] = 8'h80;
    green_mem[484] = 8'hff;
    green_mem[485] = 8'hfe;
    green_mem[486] = 8'hff;
    green_mem[487] = 8'hff;
    green_mem[488] = 8'hff;
    green_mem[489] = 8'hff;
    green_mem[490] = 8'hff;
    green_mem[491] = 8'hff;
    green_mem[492] = 8'h01;
    green_mem[493] = 8'h00;
    green_mem[494] = 8'h00;
    green_mem[495] = 8'h00;
    green_mem[496] = 8'h00;
    green_mem[497] = 8'h00;
    green_mem[498] = 8'h00;
    green_mem[499] = 8'hc0;
    green_mem[500] = 8'hff;
    green_mem[501] = 8'hff;
    green_mem[502] = 8'hff;
    green_mem[503] = 8'hff;
    green_mem[504] = 8'hff;
    green_mem[505] = 8'hff;
    green_mem[506] = 8'hff;
    green_mem[507] = 8'hff;
    green_mem[508] = 8'h03;
    green_mem[509] = 8'h00;
    green_mem[510] = 8'h00;
    green_mem[511] = 8'h00;
    green_mem[512] = 8'h00;
    green_mem[513] = 8'h00;
    green_mem[514] = 8'h00;
    green_mem[515] = 8'hc0;
    green_mem[516] = 8'hff;
    green_mem[517] = 8'hff;
    green_mem[518] = 8'hff;
    green_mem[519] = 8'hff;
    green_mem[520] = 8'hff;
    green_mem[521] = 8'hff;
    green_mem[522] = 8'hff;
    green_mem[523] = 8'hff;
    green_mem[524] = 8'h07;
    green_mem[525] = 8'h00;
    green_mem[526] = 8'h00;
    green_mem[527] = 8'h00;
    green_mem[528] = 8'h00;
    green_mem[529] = 8'h00;
    green_mem[530] = 8'h00;
    green_mem[531] = 8'hc0;
    green_mem[532] = 8'hff;
    green_mem[533] = 8'hf7;
    green_mem[534] = 8'hff;
    green_mem[535] = 8'hff;
    green_mem[536] = 8'hff;
    green_mem[537] = 8'hff;
    green_mem[538] = 8'hff;
    green_mem[539] = 8'hff;
    green_mem[540] = 8'h0f;
    green_mem[541] = 8'h00;
    green_mem[542] = 8'h00;
    green_mem[543] = 8'h00;
    green_mem[544] = 8'h00;
    green_mem[545] = 8'h00;
    green_mem[546] = 8'h00;
    green_mem[547] = 8'hf8;
    green_mem[548] = 8'hff;
    green_mem[549] = 8'hff;
    green_mem[550] = 8'hdf;
    green_mem[551] = 8'hff;
    green_mem[552] = 8'hff;
    green_mem[553] = 8'hff;
    green_mem[554] = 8'hff;
    green_mem[555] = 8'hff;
    green_mem[556] = 8'h1f;
    green_mem[557] = 8'h00;
    green_mem[558] = 8'h00;
    green_mem[559] = 8'h00;
    green_mem[560] = 8'h00;
    green_mem[561] = 8'h00;
    green_mem[562] = 8'h00;
    green_mem[563] = 8'hf8;
    green_mem[564] = 8'hff;
    green_mem[565] = 8'hff;
    green_mem[566] = 8'hfd;
    green_mem[567] = 8'hff;
    green_mem[568] = 8'hff;
    green_mem[569] = 8'hff;
    green_mem[570] = 8'hff;
    green_mem[571] = 8'hfe;
    green_mem[572] = 8'h1d;
    green_mem[573] = 8'h00;
    green_mem[574] = 8'h00;
    green_mem[575] = 8'h00;
    green_mem[576] = 8'h00;
    green_mem[577] = 8'h00;
    green_mem[578] = 8'h00;
    green_mem[579] = 8'hf0;
    green_mem[580] = 8'hff;
    green_mem[581] = 8'hff;
    green_mem[582] = 8'hff;
    green_mem[583] = 8'hff;
    green_mem[584] = 8'hff;
    green_mem[585] = 8'hff;
    green_mem[586] = 8'hff;
    green_mem[587] = 8'hff;
    green_mem[588] = 8'h7b;
    green_mem[589] = 8'h00;
    green_mem[590] = 8'h00;
    green_mem[591] = 8'h00;
    green_mem[592] = 8'h00;
    green_mem[593] = 8'h00;
    green_mem[594] = 8'h00;
    green_mem[595] = 8'hfe;
    green_mem[596] = 8'hbf;
    green_mem[597] = 8'hff;
    green_mem[598] = 8'h9f;
    green_mem[599] = 8'hff;
    green_mem[600] = 8'hff;
    green_mem[601] = 8'h0f;
    green_mem[602] = 8'hc0;
    green_mem[603] = 8'hff;
    green_mem[604] = 8'hff;
    green_mem[605] = 8'h00;
    green_mem[606] = 8'h00;
    green_mem[607] = 8'h00;
    green_mem[608] = 8'h00;
    green_mem[609] = 8'h00;
    green_mem[610] = 8'h00;
    green_mem[611] = 8'hfe;
    green_mem[612] = 8'hfd;
    green_mem[613] = 8'hff;
    green_mem[614] = 8'h07;
    green_mem[615] = 8'hff;
    green_mem[616] = 8'hff;
    green_mem[617] = 8'h00;
    green_mem[618] = 8'h00;
    green_mem[619] = 8'hfe;
    green_mem[620] = 8'hff;
    green_mem[621] = 8'h00;
    green_mem[622] = 8'h00;
    green_mem[623] = 8'h00;
    green_mem[624] = 8'h00;
    green_mem[625] = 8'h00;
    green_mem[626] = 8'h00;
    green_mem[627] = 8'hfe;
    green_mem[628] = 8'hff;
    green_mem[629] = 8'hff;
    green_mem[630] = 8'h03;
    green_mem[631] = 8'hff;
    green_mem[632] = 8'hff;
    green_mem[633] = 8'h00;
    green_mem[634] = 8'h00;
    green_mem[635] = 8'hf0;
    green_mem[636] = 8'hff;
    green_mem[637] = 8'h00;
    green_mem[638] = 8'h00;
    green_mem[639] = 8'h00;
    green_mem[640] = 8'h00;
    green_mem[641] = 8'h00;
    green_mem[642] = 8'h80;
    green_mem[643] = 8'hff;
    green_mem[644] = 8'hff;
    green_mem[645] = 8'hff;
    green_mem[646] = 8'h80;
    green_mem[647] = 8'hff;
    green_mem[648] = 8'h1f;
    green_mem[649] = 8'h00;
    green_mem[650] = 8'h00;
    green_mem[651] = 8'hf0;
    green_mem[652] = 8'hff;
    green_mem[653] = 8'h01;
    green_mem[654] = 8'h00;
    green_mem[655] = 8'h00;
    green_mem[656] = 8'h00;
    green_mem[657] = 8'h00;
    green_mem[658] = 8'h80;
    green_mem[659] = 8'hff;
    green_mem[660] = 8'hef;
    green_mem[661] = 8'hff;
    green_mem[662] = 8'h00;
    green_mem[663] = 8'hff;
    green_mem[664] = 8'h1b;
    green_mem[665] = 8'hf0;
    green_mem[666] = 8'h00;
    green_mem[667] = 8'he0;
    green_mem[668] = 8'hff;
    green_mem[669] = 8'h01;
    green_mem[670] = 8'h00;
    green_mem[671] = 8'h00;
    green_mem[672] = 8'h00;
    green_mem[673] = 8'h00;
    green_mem[674] = 8'hc0;
    green_mem[675] = 8'hff;
    green_mem[676] = 8'hef;
    green_mem[677] = 8'hfe;
    green_mem[678] = 8'h00;
    green_mem[679] = 8'hff;
    green_mem[680] = 8'h0b;
    green_mem[681] = 8'hf8;
    green_mem[682] = 8'h07;
    green_mem[683] = 8'he0;
    green_mem[684] = 8'hff;
    green_mem[685] = 8'h03;
    green_mem[686] = 8'h00;
    green_mem[687] = 8'h00;
    green_mem[688] = 8'h00;
    green_mem[689] = 8'h00;
    green_mem[690] = 8'hc0;
    green_mem[691] = 8'hbf;
    green_mem[692] = 8'hff;
    green_mem[693] = 8'h3f;
    green_mem[694] = 8'h80;
    green_mem[695] = 8'hef;
    green_mem[696] = 8'h07;
    green_mem[697] = 8'hfc;
    green_mem[698] = 8'h3f;
    green_mem[699] = 8'he0;
    green_mem[700] = 8'hff;
    green_mem[701] = 8'h07;
    green_mem[702] = 8'h00;
    green_mem[703] = 8'h00;
    green_mem[704] = 8'h00;
    green_mem[705] = 8'h00;
    green_mem[706] = 8'he0;
    green_mem[707] = 8'hff;
    green_mem[708] = 8'hff;
    green_mem[709] = 8'h3f;
    green_mem[710] = 8'ha0;
    green_mem[711] = 8'hff;
    green_mem[712] = 8'h03;
    green_mem[713] = 8'hff;
    green_mem[714] = 8'h7f;
    green_mem[715] = 8'hc0;
    green_mem[716] = 8'hff;
    green_mem[717] = 8'h07;
    green_mem[718] = 8'h00;
    green_mem[719] = 8'h00;
    green_mem[720] = 8'h00;
    green_mem[721] = 8'h00;
    green_mem[722] = 8'hc0;
    green_mem[723] = 8'hff;
    green_mem[724] = 8'hff;
    green_mem[725] = 8'h0f;
    green_mem[726] = 8'hc0;
    green_mem[727] = 8'hff;
    green_mem[728] = 8'h03;
    green_mem[729] = 8'hff;
    green_mem[730] = 8'h7f;
    green_mem[731] = 8'h88;
    green_mem[732] = 8'hff;
    green_mem[733] = 8'h0f;
    green_mem[734] = 8'h00;
    green_mem[735] = 8'h00;
    green_mem[736] = 8'h00;
    green_mem[737] = 8'h00;
    green_mem[738] = 8'hf0;
    green_mem[739] = 8'hfd;
    green_mem[740] = 8'hdf;
    green_mem[741] = 8'h0f;
    green_mem[742] = 8'h80;
    green_mem[743] = 8'hff;
    green_mem[744] = 8'h01;
    green_mem[745] = 8'hff;
    green_mem[746] = 8'hff;
    green_mem[747] = 8'h80;
    green_mem[748] = 8'hff;
    green_mem[749] = 8'h0f;
    green_mem[750] = 8'h00;
    green_mem[751] = 8'h00;
    green_mem[752] = 8'h00;
    green_mem[753] = 8'h00;
    green_mem[754] = 8'hf0;
    green_mem[755] = 8'hff;
    green_mem[756] = 8'hff;
    green_mem[757] = 8'h0f;
    green_mem[758] = 8'hc0;
    green_mem[759] = 8'hff;
    green_mem[760] = 8'h83;
    green_mem[761] = 8'hff;
    green_mem[762] = 8'hff;
    green_mem[763] = 8'h80;
    green_mem[764] = 8'hff;
    green_mem[765] = 8'h1f;
    green_mem[766] = 8'h00;
    green_mem[767] = 8'h00;
    green_mem[768] = 8'h00;
    green_mem[769] = 8'h00;
    green_mem[770] = 8'hf0;
    green_mem[771] = 8'hff;
    green_mem[772] = 8'hff;
    green_mem[773] = 8'h81;
    green_mem[774] = 8'hc0;
    green_mem[775] = 8'hff;
    green_mem[776] = 8'h01;
    green_mem[777] = 8'hff;
    green_mem[778] = 8'h7f;
    green_mem[779] = 8'h00;
    green_mem[780] = 8'hff;
    green_mem[781] = 8'h1f;
    green_mem[782] = 8'h00;
    green_mem[783] = 8'h00;
    green_mem[784] = 8'h00;
    green_mem[785] = 8'h00;
    green_mem[786] = 8'hf0;
    green_mem[787] = 8'hff;
    green_mem[788] = 8'hff;
    green_mem[789] = 8'h61;
    green_mem[790] = 8'hc0;
    green_mem[791] = 8'hff;
    green_mem[792] = 8'h01;
    green_mem[793] = 8'hfe;
    green_mem[794] = 8'hef;
    green_mem[795] = 8'h00;
    green_mem[796] = 8'hff;
    green_mem[797] = 8'h1f;
    green_mem[798] = 8'h00;
    green_mem[799] = 8'h00;
    green_mem[800] = 8'h00;
    green_mem[801] = 8'h00;
    green_mem[802] = 8'hf8;
    green_mem[803] = 8'hff;
    green_mem[804] = 8'h3f;
    green_mem[805] = 8'h70;
    green_mem[806] = 8'hc0;
    green_mem[807] = 8'hff;
    green_mem[808] = 8'h00;
    green_mem[809] = 8'hfc;
    green_mem[810] = 8'hff;
    green_mem[811] = 8'h80;
    green_mem[812] = 8'h9f;
    green_mem[813] = 8'h3f;
    green_mem[814] = 8'h00;
    green_mem[815] = 8'h00;
    green_mem[816] = 8'h00;
    green_mem[817] = 8'h00;
    green_mem[818] = 8'hfc;
    green_mem[819] = 8'hff;
    green_mem[820] = 8'h3f;
    green_mem[821] = 8'h72;
    green_mem[822] = 8'he0;
    green_mem[823] = 8'hff;
    green_mem[824] = 8'h00;
    green_mem[825] = 8'hb8;
    green_mem[826] = 8'h3f;
    green_mem[827] = 8'h00;
    green_mem[828] = 8'hff;
    green_mem[829] = 8'h3f;
    green_mem[830] = 8'h00;
    green_mem[831] = 8'h00;
    green_mem[832] = 8'h00;
    green_mem[833] = 8'h00;
    green_mem[834] = 8'hfc;
    green_mem[835] = 8'hff;
    green_mem[836] = 8'h7f;
    green_mem[837] = 8'h3c;
    green_mem[838] = 8'he0;
    green_mem[839] = 8'hfe;
    green_mem[840] = 8'h00;
    green_mem[841] = 8'hf0;
    green_mem[842] = 8'h3f;
    green_mem[843] = 8'h00;
    green_mem[844] = 8'hff;
    green_mem[845] = 8'h3f;
    green_mem[846] = 8'h00;
    green_mem[847] = 8'h00;
    green_mem[848] = 8'h00;
    green_mem[849] = 8'h00;
    green_mem[850] = 8'hfc;
    green_mem[851] = 8'hff;
    green_mem[852] = 8'h3f;
    green_mem[853] = 8'h3c;
    green_mem[854] = 8'he0;
    green_mem[855] = 8'hff;
    green_mem[856] = 8'h00;
    green_mem[857] = 8'hf8;
    green_mem[858] = 8'h3f;
    green_mem[859] = 8'h80;
    green_mem[860] = 8'hff;
    green_mem[861] = 8'h3f;
    green_mem[862] = 8'h00;
    green_mem[863] = 8'h00;
    green_mem[864] = 8'h00;
    green_mem[865] = 8'h00;
    green_mem[866] = 8'hf8;
    green_mem[867] = 8'hff;
    green_mem[868] = 8'h3f;
    green_mem[869] = 8'h7e;
    green_mem[870] = 8'he0;
    green_mem[871] = 8'hff;
    green_mem[872] = 8'h00;
    green_mem[873] = 8'hfc;
    green_mem[874] = 8'h3f;
    green_mem[875] = 8'hc4;
    green_mem[876] = 8'hff;
    green_mem[877] = 8'h3f;
    green_mem[878] = 8'h00;
    green_mem[879] = 8'h00;
    green_mem[880] = 8'h00;
    green_mem[881] = 8'h00;
    green_mem[882] = 8'hfc;
    green_mem[883] = 8'hff;
    green_mem[884] = 8'hbb;
    green_mem[885] = 8'h1f;
    green_mem[886] = 8'hf0;
    green_mem[887] = 8'hff;
    green_mem[888] = 8'h01;
    green_mem[889] = 8'hf8;
    green_mem[890] = 8'h1d;
    green_mem[891] = 8'h80;
    green_mem[892] = 8'hff;
    green_mem[893] = 8'h7f;
    green_mem[894] = 8'h00;
    green_mem[895] = 8'h00;
    green_mem[896] = 8'h00;
    green_mem[897] = 8'h00;
    green_mem[898] = 8'hfc;
    green_mem[899] = 8'hff;
    green_mem[900] = 8'hff;
    green_mem[901] = 8'h1f;
    green_mem[902] = 8'hf0;
    green_mem[903] = 8'hff;
    green_mem[904] = 8'h03;
    green_mem[905] = 8'hf8;
    green_mem[906] = 8'h1f;
    green_mem[907] = 8'hc0;
    green_mem[908] = 8'hff;
    green_mem[909] = 8'h7f;
    green_mem[910] = 8'h00;
    green_mem[911] = 8'h00;
    green_mem[912] = 8'h00;
    green_mem[913] = 8'h00;
    green_mem[914] = 8'hfe;
    green_mem[915] = 8'hff;
    green_mem[916] = 8'hff;
    green_mem[917] = 8'h1f;
    green_mem[918] = 8'he0;
    green_mem[919] = 8'hff;
    green_mem[920] = 8'h03;
    green_mem[921] = 8'hfe;
    green_mem[922] = 8'h0f;
    green_mem[923] = 8'hf0;
    green_mem[924] = 8'hff;
    green_mem[925] = 8'h7f;
    green_mem[926] = 8'h00;
    green_mem[927] = 8'h00;
    green_mem[928] = 8'h00;
    green_mem[929] = 8'h00;
    green_mem[930] = 8'hfc;
    green_mem[931] = 8'hff;
    green_mem[932] = 8'hff;
    green_mem[933] = 8'h1f;
    green_mem[934] = 8'hf0;
    green_mem[935] = 8'hff;
    green_mem[936] = 8'h9f;
    green_mem[937] = 8'hff;
    green_mem[938] = 8'h07;
    green_mem[939] = 8'hf0;
    green_mem[940] = 8'hff;
    green_mem[941] = 8'h7f;
    green_mem[942] = 8'h00;
    green_mem[943] = 8'h00;
    green_mem[944] = 8'h00;
    green_mem[945] = 8'h00;
    green_mem[946] = 8'hfc;
    green_mem[947] = 8'hff;
    green_mem[948] = 8'hff;
    green_mem[949] = 8'h0f;
    green_mem[950] = 8'hf0;
    green_mem[951] = 8'hff;
    green_mem[952] = 8'hff;
    green_mem[953] = 8'h7f;
    green_mem[954] = 8'h01;
    green_mem[955] = 8'hf8;
    green_mem[956] = 8'hff;
    green_mem[957] = 8'hff;
    green_mem[958] = 8'h00;
    green_mem[959] = 8'h00;
    green_mem[960] = 8'h00;
    green_mem[961] = 8'h00;
    green_mem[962] = 8'hf0;
    green_mem[963] = 8'hff;
    green_mem[964] = 8'hff;
    green_mem[965] = 8'h87;
    green_mem[966] = 8'hf8;
    green_mem[967] = 8'hff;
    green_mem[968] = 8'hff;
    green_mem[969] = 8'h7f;
    green_mem[970] = 8'h00;
    green_mem[971] = 8'hfc;
    green_mem[972] = 8'hff;
    green_mem[973] = 8'hff;
    green_mem[974] = 8'h00;
    green_mem[975] = 8'h00;
    green_mem[976] = 8'h00;
    green_mem[977] = 8'h00;
    green_mem[978] = 8'hff;
    green_mem[979] = 8'hff;
    green_mem[980] = 8'hff;
    green_mem[981] = 8'h0f;
    green_mem[982] = 8'hf8;
    green_mem[983] = 8'hff;
    green_mem[984] = 8'hff;
    green_mem[985] = 8'h77;
    green_mem[986] = 8'h00;
    green_mem[987] = 8'hff;
    green_mem[988] = 8'hfd;
    green_mem[989] = 8'h7f;
    green_mem[990] = 8'h00;
    green_mem[991] = 8'h00;
    green_mem[992] = 8'h00;
    green_mem[993] = 8'h00;
    green_mem[994] = 8'hff;
    green_mem[995] = 8'hff;
    green_mem[996] = 8'hff;
    green_mem[997] = 8'h0f;
    green_mem[998] = 8'hf8;
    green_mem[999] = 8'hff;
    green_mem[1000] = 8'hff;
    green_mem[1001] = 8'h7f;
    green_mem[1002] = 8'h00;
    green_mem[1003] = 8'hff;
    green_mem[1004] = 8'hef;
    green_mem[1005] = 8'h7f;
    green_mem[1006] = 8'h00;
    green_mem[1007] = 8'h00;
    green_mem[1008] = 8'h00;
    green_mem[1009] = 8'h00;
    green_mem[1010] = 8'hff;
    green_mem[1011] = 8'hff;
    green_mem[1012] = 8'hff;
    green_mem[1013] = 8'h0f;
    green_mem[1014] = 8'hf8;
    green_mem[1015] = 8'hff;
    green_mem[1016] = 8'hff;
    green_mem[1017] = 8'h1f;
    green_mem[1018] = 8'he0;
    green_mem[1019] = 8'hff;
    green_mem[1020] = 8'hff;
    green_mem[1021] = 8'h3f;
    green_mem[1022] = 8'h00;
    green_mem[1023] = 8'h00;
    green_mem[1024] = 8'h00;
    green_mem[1025] = 8'h00;
    green_mem[1026] = 8'hfe;
    green_mem[1027] = 8'hff;
    green_mem[1028] = 8'hff;
    green_mem[1029] = 8'h07;
    green_mem[1030] = 8'h7c;
    green_mem[1031] = 8'hff;
    green_mem[1032] = 8'hff;
    green_mem[1033] = 8'h0f;
    green_mem[1034] = 8'hf0;
    green_mem[1035] = 8'hff;
    green_mem[1036] = 8'hff;
    green_mem[1037] = 8'h7f;
    green_mem[1038] = 8'h00;
    green_mem[1039] = 8'h00;
    green_mem[1040] = 8'h00;
    green_mem[1041] = 8'h00;
    green_mem[1042] = 8'hfe;
    green_mem[1043] = 8'hff;
    green_mem[1044] = 8'hff;
    green_mem[1045] = 8'h07;
    green_mem[1046] = 8'hf8;
    green_mem[1047] = 8'hff;
    green_mem[1048] = 8'hff;
    green_mem[1049] = 8'h03;
    green_mem[1050] = 8'hf6;
    green_mem[1051] = 8'hff;
    green_mem[1052] = 8'hff;
    green_mem[1053] = 8'he7;
    green_mem[1054] = 8'h00;
    green_mem[1055] = 8'h00;
    green_mem[1056] = 8'h00;
    green_mem[1057] = 8'h00;
    green_mem[1058] = 8'hfe;
    green_mem[1059] = 8'hff;
    green_mem[1060] = 8'hff;
    green_mem[1061] = 8'h47;
    green_mem[1062] = 8'hfc;
    green_mem[1063] = 8'hff;
    green_mem[1064] = 8'hff;
    green_mem[1065] = 8'h43;
    green_mem[1066] = 8'hff;
    green_mem[1067] = 8'hff;
    green_mem[1068] = 8'hff;
    green_mem[1069] = 8'h7f;
    green_mem[1070] = 8'h00;
    green_mem[1071] = 8'h00;
    green_mem[1072] = 8'h00;
    green_mem[1073] = 8'h00;
    green_mem[1074] = 8'hfe;
    green_mem[1075] = 8'hbf;
    green_mem[1076] = 8'hff;
    green_mem[1077] = 8'h03;
    green_mem[1078] = 8'hfe;
    green_mem[1079] = 8'hff;
    green_mem[1080] = 8'h7e;
    green_mem[1081] = 8'he0;
    green_mem[1082] = 8'hff;
    green_mem[1083] = 8'hff;
    green_mem[1084] = 8'hff;
    green_mem[1085] = 8'h7f;
    green_mem[1086] = 8'h00;
    green_mem[1087] = 8'h00;
    green_mem[1088] = 8'h00;
    green_mem[1089] = 8'h00;
    green_mem[1090] = 8'hfe;
    green_mem[1091] = 8'hff;
    green_mem[1092] = 8'hff;
    green_mem[1093] = 8'h03;
    green_mem[1094] = 8'hfe;
    green_mem[1095] = 8'hff;
    green_mem[1096] = 8'h7e;
    green_mem[1097] = 8'he0;
    green_mem[1098] = 8'hef;
    green_mem[1099] = 8'hff;
    green_mem[1100] = 8'hff;
    green_mem[1101] = 8'hff;
    green_mem[1102] = 8'h00;
    green_mem[1103] = 8'h00;
    green_mem[1104] = 8'h00;
    green_mem[1105] = 8'h00;
    green_mem[1106] = 8'hfc;
    green_mem[1107] = 8'hff;
    green_mem[1108] = 8'hf7;
    green_mem[1109] = 8'h03;
    green_mem[1110] = 8'hfe;
    green_mem[1111] = 8'hff;
    green_mem[1112] = 8'h1f;
    green_mem[1113] = 8'h7c;
    green_mem[1114] = 8'hff;
    green_mem[1115] = 8'hff;
    green_mem[1116] = 8'hff;
    green_mem[1117] = 8'h7f;
    green_mem[1118] = 8'h00;
    green_mem[1119] = 8'h00;
    green_mem[1120] = 8'h00;
    green_mem[1121] = 8'h00;
    green_mem[1122] = 8'hfc;
    green_mem[1123] = 8'hbf;
    green_mem[1124] = 8'hff;
    green_mem[1125] = 8'h83;
    green_mem[1126] = 8'hff;
    green_mem[1127] = 8'hff;
    green_mem[1128] = 8'h07;
    green_mem[1129] = 8'hfc;
    green_mem[1130] = 8'hff;
    green_mem[1131] = 8'hff;
    green_mem[1132] = 8'hff;
    green_mem[1133] = 8'h7f;
    green_mem[1134] = 8'h00;
    green_mem[1135] = 8'h00;
    green_mem[1136] = 8'h00;
    green_mem[1137] = 8'h00;
    green_mem[1138] = 8'hfe;
    green_mem[1139] = 8'hff;
    green_mem[1140] = 8'hff;
    green_mem[1141] = 8'h03;
    green_mem[1142] = 8'hfe;
    green_mem[1143] = 8'hff;
    green_mem[1144] = 8'h87;
    green_mem[1145] = 8'hff;
    green_mem[1146] = 8'hff;
    green_mem[1147] = 8'hff;
    green_mem[1148] = 8'hff;
    green_mem[1149] = 8'h7f;
    green_mem[1150] = 8'h00;
    green_mem[1151] = 8'h00;
    green_mem[1152] = 8'h00;
    green_mem[1153] = 8'h00;
    green_mem[1154] = 8'hfe;
    green_mem[1155] = 8'hff;
    green_mem[1156] = 8'hff;
    green_mem[1157] = 8'h03;
    green_mem[1158] = 8'hfe;
    green_mem[1159] = 8'hfb;
    green_mem[1160] = 8'h80;
    green_mem[1161] = 8'hff;
    green_mem[1162] = 8'hff;
    green_mem[1163] = 8'hff;
    green_mem[1164] = 8'hff;
    green_mem[1165] = 8'h7f;
    green_mem[1166] = 8'h00;
    green_mem[1167] = 8'h00;
    green_mem[1168] = 8'h00;
    green_mem[1169] = 8'h00;
    green_mem[1170] = 8'hfc;
    green_mem[1171] = 8'hff;
    green_mem[1172] = 8'hff;
    green_mem[1173] = 8'h03;
    green_mem[1174] = 8'hfe;
    green_mem[1175] = 8'h7f;
    green_mem[1176] = 8'h80;
    green_mem[1177] = 8'hfd;
    green_mem[1178] = 8'hef;
    green_mem[1179] = 8'hff;
    green_mem[1180] = 8'hff;
    green_mem[1181] = 8'h7e;
    green_mem[1182] = 8'h00;
    green_mem[1183] = 8'h00;
    green_mem[1184] = 8'h00;
    green_mem[1185] = 8'h00;
    green_mem[1186] = 8'hfc;
    green_mem[1187] = 8'hff;
    green_mem[1188] = 8'hff;
    green_mem[1189] = 8'h03;
    green_mem[1190] = 8'hfe;
    green_mem[1191] = 8'h7f;
    green_mem[1192] = 8'h00;
    green_mem[1193] = 8'hf8;
    green_mem[1194] = 8'hef;
    green_mem[1195] = 8'hc7;
    green_mem[1196] = 8'hff;
    green_mem[1197] = 8'h3f;
    green_mem[1198] = 8'h00;
    green_mem[1199] = 8'h00;
    green_mem[1200] = 8'h00;
    green_mem[1201] = 8'h00;
    green_mem[1202] = 8'hf8;
    green_mem[1203] = 8'h7f;
    green_mem[1204] = 8'hcf;
    green_mem[1205] = 8'h03;
    green_mem[1206] = 8'hfe;
    green_mem[1207] = 8'h7f;
    green_mem[1208] = 8'h00;
    green_mem[1209] = 8'h80;
    green_mem[1210] = 8'hff;
    green_mem[1211] = 8'hc3;
    green_mem[1212] = 8'hff;
    green_mem[1213] = 8'h37;
    green_mem[1214] = 8'h00;
    green_mem[1215] = 8'h00;
    green_mem[1216] = 8'h00;
    green_mem[1217] = 8'h00;
    green_mem[1218] = 8'hf8;
    green_mem[1219] = 8'hff;
    green_mem[1220] = 8'hff;
    green_mem[1221] = 8'h01;
    green_mem[1222] = 8'hff;
    green_mem[1223] = 8'h0f;
    green_mem[1224] = 8'h00;
    green_mem[1225] = 8'h00;
    green_mem[1226] = 8'hf8;
    green_mem[1227] = 8'hf1;
    green_mem[1228] = 8'hff;
    green_mem[1229] = 8'h3f;
    green_mem[1230] = 8'h00;
    green_mem[1231] = 8'h00;
    green_mem[1232] = 8'h00;
    green_mem[1233] = 8'h00;
    green_mem[1234] = 8'hb8;
    green_mem[1235] = 8'hff;
    green_mem[1236] = 8'hff;
    green_mem[1237] = 8'h80;
    green_mem[1238] = 8'hff;
    green_mem[1239] = 8'h07;
    green_mem[1240] = 8'h08;
    green_mem[1241] = 8'h00;
    green_mem[1242] = 8'h38;
    green_mem[1243] = 8'hf0;
    green_mem[1244] = 8'hff;
    green_mem[1245] = 8'h1f;
    green_mem[1246] = 8'h00;
    green_mem[1247] = 8'h00;
    green_mem[1248] = 8'h00;
    green_mem[1249] = 8'h00;
    green_mem[1250] = 8'hf0;
    green_mem[1251] = 8'hdf;
    green_mem[1252] = 8'hff;
    green_mem[1253] = 8'h90;
    green_mem[1254] = 8'hff;
    green_mem[1255] = 8'h07;
    green_mem[1256] = 8'h00;
    green_mem[1257] = 8'h00;
    green_mem[1258] = 8'h00;
    green_mem[1259] = 8'hf8;
    green_mem[1260] = 8'hef;
    green_mem[1261] = 8'h1f;
    green_mem[1262] = 8'h00;
    green_mem[1263] = 8'h00;
    green_mem[1264] = 8'h00;
    green_mem[1265] = 8'h00;
    green_mem[1266] = 8'hf0;
    green_mem[1267] = 8'hff;
    green_mem[1268] = 8'hff;
    green_mem[1269] = 8'hc0;
    green_mem[1270] = 8'hff;
    green_mem[1271] = 8'h07;
    green_mem[1272] = 8'h00;
    green_mem[1273] = 8'h00;
    green_mem[1274] = 8'h00;
    green_mem[1275] = 8'hf8;
    green_mem[1276] = 8'hff;
    green_mem[1277] = 8'h1f;
    green_mem[1278] = 8'h00;
    green_mem[1279] = 8'h00;
    green_mem[1280] = 8'h00;
    green_mem[1281] = 8'h00;
    green_mem[1282] = 8'hf0;
    green_mem[1283] = 8'hff;
    green_mem[1284] = 8'hff;
    green_mem[1285] = 8'h80;
    green_mem[1286] = 8'hff;
    green_mem[1287] = 8'h03;
    green_mem[1288] = 8'h18;
    green_mem[1289] = 8'h00;
    green_mem[1290] = 8'h00;
    green_mem[1291] = 8'hfc;
    green_mem[1292] = 8'hff;
    green_mem[1293] = 8'h0f;
    green_mem[1294] = 8'h00;
    green_mem[1295] = 8'h00;
    green_mem[1296] = 8'h00;
    green_mem[1297] = 8'h00;
    green_mem[1298] = 8'he0;
    green_mem[1299] = 8'hff;
    green_mem[1300] = 8'h37;
    green_mem[1301] = 8'h00;
    green_mem[1302] = 8'hff;
    green_mem[1303] = 8'h80;
    green_mem[1304] = 8'hff;
    green_mem[1305] = 8'h00;
    green_mem[1306] = 8'h00;
    green_mem[1307] = 8'hfc;
    green_mem[1308] = 8'hff;
    green_mem[1309] = 8'h0f;
    green_mem[1310] = 8'h00;
    green_mem[1311] = 8'h00;
    green_mem[1312] = 8'h00;
    green_mem[1313] = 8'h00;
    green_mem[1314] = 8'he0;
    green_mem[1315] = 8'hff;
    green_mem[1316] = 8'h03;
    green_mem[1317] = 8'h00;
    green_mem[1318] = 8'hf0;
    green_mem[1319] = 8'hf0;
    green_mem[1320] = 8'hff;
    green_mem[1321] = 8'h03;
    green_mem[1322] = 8'h80;
    green_mem[1323] = 8'hff;
    green_mem[1324] = 8'hdf;
    green_mem[1325] = 8'h0f;
    green_mem[1326] = 8'h00;
    green_mem[1327] = 8'h00;
    green_mem[1328] = 8'h00;
    green_mem[1329] = 8'h00;
    green_mem[1330] = 8'he0;
    green_mem[1331] = 8'hff;
    green_mem[1332] = 8'h03;
    green_mem[1333] = 8'h00;
    green_mem[1334] = 8'hf0;
    green_mem[1335] = 8'hf8;
    green_mem[1336] = 8'hff;
    green_mem[1337] = 8'h0f;
    green_mem[1338] = 8'hc0;
    green_mem[1339] = 8'hff;
    green_mem[1340] = 8'hff;
    green_mem[1341] = 8'h07;
    green_mem[1342] = 8'h00;
    green_mem[1343] = 8'h00;
    green_mem[1344] = 8'h00;
    green_mem[1345] = 8'h00;
    green_mem[1346] = 8'h80;
    green_mem[1347] = 8'hff;
    green_mem[1348] = 8'h43;
    green_mem[1349] = 8'h86;
    green_mem[1350] = 8'hf8;
    green_mem[1351] = 8'hfd;
    green_mem[1352] = 8'hff;
    green_mem[1353] = 8'hff;
    green_mem[1354] = 8'hfb;
    green_mem[1355] = 8'hff;
    green_mem[1356] = 8'hff;
    green_mem[1357] = 8'h07;
    green_mem[1358] = 8'h00;
    green_mem[1359] = 8'h00;
    green_mem[1360] = 8'h00;
    green_mem[1361] = 8'h00;
    green_mem[1362] = 8'h80;
    green_mem[1363] = 8'hff;
    green_mem[1364] = 8'hf7;
    green_mem[1365] = 8'hc7;
    green_mem[1366] = 8'hfd;
    green_mem[1367] = 8'hff;
    green_mem[1368] = 8'hff;
    green_mem[1369] = 8'hff;
    green_mem[1370] = 8'hff;
    green_mem[1371] = 8'hff;
    green_mem[1372] = 8'hff;
    green_mem[1373] = 8'h07;
    green_mem[1374] = 8'h00;
    green_mem[1375] = 8'h00;
    green_mem[1376] = 8'h00;
    green_mem[1377] = 8'h00;
    green_mem[1378] = 8'hc0;
    green_mem[1379] = 8'hff;
    green_mem[1380] = 8'hff;
    green_mem[1381] = 8'hff;
    green_mem[1382] = 8'hfd;
    green_mem[1383] = 8'hf7;
    green_mem[1384] = 8'hff;
    green_mem[1385] = 8'hff;
    green_mem[1386] = 8'hff;
    green_mem[1387] = 8'hff;
    green_mem[1388] = 8'hff;
    green_mem[1389] = 8'h07;
    green_mem[1390] = 8'h00;
    green_mem[1391] = 8'h00;
    green_mem[1392] = 8'h00;
    green_mem[1393] = 8'h00;
    green_mem[1394] = 8'h00;
    green_mem[1395] = 8'hff;
    green_mem[1396] = 8'hff;
    green_mem[1397] = 8'hfd;
    green_mem[1398] = 8'hff;
    green_mem[1399] = 8'hf7;
    green_mem[1400] = 8'hff;
    green_mem[1401] = 8'hff;
    green_mem[1402] = 8'hff;
    green_mem[1403] = 8'hff;
    green_mem[1404] = 8'hff;
    green_mem[1405] = 8'h03;
    green_mem[1406] = 8'h00;
    green_mem[1407] = 8'h00;
    green_mem[1408] = 8'h00;
    green_mem[1409] = 8'h00;
    green_mem[1410] = 8'h00;
    green_mem[1411] = 8'hff;
    green_mem[1412] = 8'hff;
    green_mem[1413] = 8'hff;
    green_mem[1414] = 8'hff;
    green_mem[1415] = 8'hff;
    green_mem[1416] = 8'hff;
    green_mem[1417] = 8'hff;
    green_mem[1418] = 8'hf7;
    green_mem[1419] = 8'hff;
    green_mem[1420] = 8'hff;
    green_mem[1421] = 8'h00;
    green_mem[1422] = 8'h00;
    green_mem[1423] = 8'h00;
    green_mem[1424] = 8'h00;
    green_mem[1425] = 8'h00;
    green_mem[1426] = 8'h00;
    green_mem[1427] = 8'hff;
    green_mem[1428] = 8'hfe;
    green_mem[1429] = 8'hf7;
    green_mem[1430] = 8'hff;
    green_mem[1431] = 8'hff;
    green_mem[1432] = 8'hff;
    green_mem[1433] = 8'hff;
    green_mem[1434] = 8'hff;
    green_mem[1435] = 8'hff;
    green_mem[1436] = 8'hff;
    green_mem[1437] = 8'h00;
    green_mem[1438] = 8'h00;
    green_mem[1439] = 8'h00;
    green_mem[1440] = 8'h00;
    green_mem[1441] = 8'h00;
    green_mem[1442] = 8'h00;
    green_mem[1443] = 8'hfc;
    green_mem[1444] = 8'hef;
    green_mem[1445] = 8'hff;
    green_mem[1446] = 8'hff;
    green_mem[1447] = 8'hff;
    green_mem[1448] = 8'hff;
    green_mem[1449] = 8'hff;
    green_mem[1450] = 8'hff;
    green_mem[1451] = 8'hff;
    green_mem[1452] = 8'hff;
    green_mem[1453] = 8'h00;
    green_mem[1454] = 8'h00;
    green_mem[1455] = 8'h00;
    green_mem[1456] = 8'h00;
    green_mem[1457] = 8'h00;
    green_mem[1458] = 8'h00;
    green_mem[1459] = 8'hfc;
    green_mem[1460] = 8'hff;
    green_mem[1461] = 8'hff;
    green_mem[1462] = 8'hff;
    green_mem[1463] = 8'hff;
    green_mem[1464] = 8'h9f;
    green_mem[1465] = 8'hff;
    green_mem[1466] = 8'hff;
    green_mem[1467] = 8'hff;
    green_mem[1468] = 8'h3f;
    green_mem[1469] = 8'h00;
    green_mem[1470] = 8'h00;
    green_mem[1471] = 8'h00;
    green_mem[1472] = 8'h00;
    green_mem[1473] = 8'h00;
    green_mem[1474] = 8'h00;
    green_mem[1475] = 8'hf8;
    green_mem[1476] = 8'hff;
    green_mem[1477] = 8'hff;
    green_mem[1478] = 8'hff;
    green_mem[1479] = 8'hff;
    green_mem[1480] = 8'hff;
    green_mem[1481] = 8'hff;
    green_mem[1482] = 8'hff;
    green_mem[1483] = 8'hff;
    green_mem[1484] = 8'h3f;
    green_mem[1485] = 8'h00;
    green_mem[1486] = 8'h00;
    green_mem[1487] = 8'h00;
    green_mem[1488] = 8'h00;
    green_mem[1489] = 8'h00;
    green_mem[1490] = 8'h00;
    green_mem[1491] = 8'h70;
    green_mem[1492] = 8'h7f;
    green_mem[1493] = 8'hff;
    green_mem[1494] = 8'hff;
    green_mem[1495] = 8'hff;
    green_mem[1496] = 8'hf7;
    green_mem[1497] = 8'hff;
    green_mem[1498] = 8'hff;
    green_mem[1499] = 8'hf7;
    green_mem[1500] = 8'h1f;
    green_mem[1501] = 8'h00;
    green_mem[1502] = 8'h00;
    green_mem[1503] = 8'h00;
    green_mem[1504] = 8'h00;
    green_mem[1505] = 8'h00;
    green_mem[1506] = 8'h00;
    green_mem[1507] = 8'he0;
    green_mem[1508] = 8'hff;
    green_mem[1509] = 8'hff;
    green_mem[1510] = 8'hff;
    green_mem[1511] = 8'hff;
    green_mem[1512] = 8'hf7;
    green_mem[1513] = 8'hef;
    green_mem[1514] = 8'hff;
    green_mem[1515] = 8'hff;
    green_mem[1516] = 8'h0f;
    green_mem[1517] = 8'h00;
    green_mem[1518] = 8'h00;
    green_mem[1519] = 8'h00;
    green_mem[1520] = 8'h00;
    green_mem[1521] = 8'h00;
    green_mem[1522] = 8'h00;
    green_mem[1523] = 8'he0;
    green_mem[1524] = 8'hfd;
    green_mem[1525] = 8'hff;
    green_mem[1526] = 8'hff;
    green_mem[1527] = 8'hff;
    green_mem[1528] = 8'hff;
    green_mem[1529] = 8'hff;
    green_mem[1530] = 8'hff;
    green_mem[1531] = 8'hff;
    green_mem[1532] = 8'h03;
    green_mem[1533] = 8'h00;
    green_mem[1534] = 8'h00;
    green_mem[1535] = 8'h00;
    green_mem[1536] = 8'h00;
    green_mem[1537] = 8'h00;
    green_mem[1538] = 8'h00;
    green_mem[1539] = 8'hc0;
    green_mem[1540] = 8'hff;
    green_mem[1541] = 8'hff;
    green_mem[1542] = 8'hff;
    green_mem[1543] = 8'hef;
    green_mem[1544] = 8'hff;
    green_mem[1545] = 8'hff;
    green_mem[1546] = 8'h7b;
    green_mem[1547] = 8'hff;
    green_mem[1548] = 8'h01;
    green_mem[1549] = 8'h00;
    green_mem[1550] = 8'h00;
    green_mem[1551] = 8'h00;
    green_mem[1552] = 8'h00;
    green_mem[1553] = 8'h00;
    green_mem[1554] = 8'h00;
    green_mem[1555] = 8'h00;
    green_mem[1556] = 8'hff;
    green_mem[1557] = 8'hff;
    green_mem[1558] = 8'hff;
    green_mem[1559] = 8'hff;
    green_mem[1560] = 8'hff;
    green_mem[1561] = 8'hff;
    green_mem[1562] = 8'hff;
    green_mem[1563] = 8'hff;
    green_mem[1564] = 8'h00;
    green_mem[1565] = 8'h00;
    green_mem[1566] = 8'h00;
    green_mem[1567] = 8'h00;
    green_mem[1568] = 8'h00;
    green_mem[1569] = 8'h00;
    green_mem[1570] = 8'h00;
    green_mem[1571] = 8'h00;
    green_mem[1572] = 8'hef;
    green_mem[1573] = 8'hff;
    green_mem[1574] = 8'hff;
    green_mem[1575] = 8'hff;
    green_mem[1576] = 8'hff;
    green_mem[1577] = 8'hff;
    green_mem[1578] = 8'hff;
    green_mem[1579] = 8'hff;
    green_mem[1580] = 8'h00;
    green_mem[1581] = 8'h00;
    green_mem[1582] = 8'h00;
    green_mem[1583] = 8'h00;
    green_mem[1584] = 8'h00;
    green_mem[1585] = 8'h00;
    green_mem[1586] = 8'h00;
    green_mem[1587] = 8'h00;
    green_mem[1588] = 8'hfe;
    green_mem[1589] = 8'hff;
    green_mem[1590] = 8'hff;
    green_mem[1591] = 8'hff;
    green_mem[1592] = 8'hff;
    green_mem[1593] = 8'hff;
    green_mem[1594] = 8'hff;
    green_mem[1595] = 8'h7f;
    green_mem[1596] = 8'h00;
    green_mem[1597] = 8'h00;
    green_mem[1598] = 8'h00;
    green_mem[1599] = 8'h00;
    green_mem[1600] = 8'h00;
    green_mem[1601] = 8'h00;
    green_mem[1602] = 8'h00;
    green_mem[1603] = 8'h00;
    green_mem[1604] = 8'hf0;
    green_mem[1605] = 8'hff;
    green_mem[1606] = 8'hff;
    green_mem[1607] = 8'hff;
    green_mem[1608] = 8'hff;
    green_mem[1609] = 8'hff;
    green_mem[1610] = 8'hff;
    green_mem[1611] = 8'h1f;
    green_mem[1612] = 8'h00;
    green_mem[1613] = 8'h00;
    green_mem[1614] = 8'h00;
    green_mem[1615] = 8'h00;
    green_mem[1616] = 8'h00;
    green_mem[1617] = 8'h00;
    green_mem[1618] = 8'h00;
    green_mem[1619] = 8'h00;
    green_mem[1620] = 8'hf0;
    green_mem[1621] = 8'hff;
    green_mem[1622] = 8'hff;
    green_mem[1623] = 8'hff;
    green_mem[1624] = 8'hf7;
    green_mem[1625] = 8'hff;
    green_mem[1626] = 8'hff;
    green_mem[1627] = 8'h1f;
    green_mem[1628] = 8'h00;
    green_mem[1629] = 8'h00;
    green_mem[1630] = 8'h00;
    green_mem[1631] = 8'h00;
    green_mem[1632] = 8'h00;
    green_mem[1633] = 8'h00;
    green_mem[1634] = 8'h00;
    green_mem[1635] = 8'h00;
    green_mem[1636] = 8'he0;
    green_mem[1637] = 8'hff;
    green_mem[1638] = 8'hf6;
    green_mem[1639] = 8'hef;
    green_mem[1640] = 8'hff;
    green_mem[1641] = 8'hfd;
    green_mem[1642] = 8'hff;
    green_mem[1643] = 8'h07;
    green_mem[1644] = 8'h00;
    green_mem[1645] = 8'h00;
    green_mem[1646] = 8'h00;
    green_mem[1647] = 8'h00;
    green_mem[1648] = 8'h00;
    green_mem[1649] = 8'h00;
    green_mem[1650] = 8'h00;
    green_mem[1651] = 8'h00;
    green_mem[1652] = 8'h00;
    green_mem[1653] = 8'h7e;
    green_mem[1654] = 8'hff;
    green_mem[1655] = 8'hff;
    green_mem[1656] = 8'hff;
    green_mem[1657] = 8'hff;
    green_mem[1658] = 8'hff;
    green_mem[1659] = 8'h03;
    green_mem[1660] = 8'h00;
    green_mem[1661] = 8'h00;
    green_mem[1662] = 8'h00;
    green_mem[1663] = 8'h00;
    green_mem[1664] = 8'h00;
    green_mem[1665] = 8'h00;
    green_mem[1666] = 8'h00;
    green_mem[1667] = 8'h00;
    green_mem[1668] = 8'h00;
    green_mem[1669] = 8'hfe;
    green_mem[1670] = 8'hff;
    green_mem[1671] = 8'hff;
    green_mem[1672] = 8'hcf;
    green_mem[1673] = 8'hff;
    green_mem[1674] = 8'hff;
    green_mem[1675] = 8'h00;
    green_mem[1676] = 8'h00;
    green_mem[1677] = 8'h00;
    green_mem[1678] = 8'h00;
    green_mem[1679] = 8'h00;
    green_mem[1680] = 8'h00;
    green_mem[1681] = 8'h00;
    green_mem[1682] = 8'h00;
    green_mem[1683] = 8'h00;
    green_mem[1684] = 8'h00;
    green_mem[1685] = 8'hf8;
    green_mem[1686] = 8'hff;
    green_mem[1687] = 8'hdf;
    green_mem[1688] = 8'hff;
    green_mem[1689] = 8'hfc;
    green_mem[1690] = 8'h3f;
    green_mem[1691] = 8'h00;
    green_mem[1692] = 8'h00;
    green_mem[1693] = 8'h00;
    green_mem[1694] = 8'h00;
    green_mem[1695] = 8'h00;
    green_mem[1696] = 8'h00;
    green_mem[1697] = 8'h00;
    green_mem[1698] = 8'h00;
    green_mem[1699] = 8'h00;
    green_mem[1700] = 8'h00;
    green_mem[1701] = 8'hf0;
    green_mem[1702] = 8'hff;
    green_mem[1703] = 8'hff;
    green_mem[1704] = 8'hfb;
    green_mem[1705] = 8'hff;
    green_mem[1706] = 8'h1f;
    green_mem[1707] = 8'h00;
    green_mem[1708] = 8'h00;
    green_mem[1709] = 8'h00;
    green_mem[1710] = 8'h00;
    green_mem[1711] = 8'h00;
    green_mem[1712] = 8'h00;
    green_mem[1713] = 8'h00;
    green_mem[1714] = 8'h00;
    green_mem[1715] = 8'h00;
    green_mem[1716] = 8'h00;
    green_mem[1717] = 8'h00;
    green_mem[1718] = 8'hff;
    green_mem[1719] = 8'hff;
    green_mem[1720] = 8'hff;
    green_mem[1721] = 8'hff;
    green_mem[1722] = 8'h01;
    green_mem[1723] = 8'h00;
    green_mem[1724] = 8'h00;
    green_mem[1725] = 8'h00;
    green_mem[1726] = 8'h00;
    green_mem[1727] = 8'h00;
    green_mem[1728] = 8'h00;
    green_mem[1729] = 8'h00;
    green_mem[1730] = 8'h00;
    green_mem[1731] = 8'h00;
    green_mem[1732] = 8'h00;
    green_mem[1733] = 8'h00;
    green_mem[1734] = 8'hfe;
    green_mem[1735] = 8'hff;
    green_mem[1736] = 8'hff;
    green_mem[1737] = 8'h3f;
    green_mem[1738] = 8'h00;
    green_mem[1739] = 8'h00;
    green_mem[1740] = 8'h00;
    green_mem[1741] = 8'h00;
    green_mem[1742] = 8'h00;
    green_mem[1743] = 8'h00;
    green_mem[1744] = 8'h00;
    green_mem[1745] = 8'h00;
    green_mem[1746] = 8'h00;
    green_mem[1747] = 8'h00;
    green_mem[1748] = 8'h00;
    green_mem[1749] = 8'h00;
    green_mem[1750] = 8'h18;
    green_mem[1751] = 8'hfe;
    green_mem[1752] = 8'hff;
    green_mem[1753] = 8'h1f;
    green_mem[1754] = 8'h00;
    green_mem[1755] = 8'h00;
    green_mem[1756] = 8'h00;
    green_mem[1757] = 8'h00;
    green_mem[1758] = 8'h00;
    green_mem[1759] = 8'h00;
    green_mem[1760] = 8'h00;
    green_mem[1761] = 8'h00;
    green_mem[1762] = 8'h00;
    green_mem[1763] = 8'h00;
    green_mem[1764] = 8'h00;
    green_mem[1765] = 8'h00;
    green_mem[1766] = 8'h00;
    green_mem[1767] = 8'hee;
    green_mem[1768] = 8'hff;
    green_mem[1769] = 8'h00;
    green_mem[1770] = 8'h00;
    green_mem[1771] = 8'h00;
    green_mem[1772] = 8'h00;
    green_mem[1773] = 8'h00;
    green_mem[1774] = 8'h00;
    green_mem[1775] = 8'h00;
    green_mem[1776] = 8'h00;
    green_mem[1777] = 8'h00;
    green_mem[1778] = 8'h00;
    green_mem[1779] = 8'h00;
    green_mem[1780] = 8'h00;
    green_mem[1781] = 8'h00;
    green_mem[1782] = 8'h00;
    green_mem[1783] = 8'h00;
    green_mem[1784] = 8'h0c;
    green_mem[1785] = 8'h00;
    green_mem[1786] = 8'h00;
    green_mem[1787] = 8'h00;
    green_mem[1788] = 8'h00;
    green_mem[1789] = 8'h00;
    green_mem[1790] = 8'h00;
    green_mem[1791] = 8'h00;
    green_mem[1792] = 8'h00;
    green_mem[1793] = 8'h00;
    green_mem[1794] = 8'h00;
    green_mem[1795] = 8'h00;
    green_mem[1796] = 8'h00;
    green_mem[1797] = 8'h00;
    green_mem[1798] = 8'h00;
    green_mem[1799] = 8'h00;
    green_mem[1800] = 8'h00;
    green_mem[1801] = 8'h00;
    green_mem[1802] = 8'h00;
    green_mem[1803] = 8'h00;
    green_mem[1804] = 8'h00;
    green_mem[1805] = 8'h00;
    green_mem[1806] = 8'h00;
    green_mem[1807] = 8'h00;
    green_mem[1808] = 8'h00;
    green_mem[1809] = 8'h00;
    green_mem[1810] = 8'h00;
    green_mem[1811] = 8'h00;
    green_mem[1812] = 8'h00;
    green_mem[1813] = 8'h00;
    green_mem[1814] = 8'h00;
    green_mem[1815] = 8'h00;
    green_mem[1816] = 8'h00;
    green_mem[1817] = 8'h00;
    green_mem[1818] = 8'h00;
    green_mem[1819] = 8'h00;
    green_mem[1820] = 8'h00;
    green_mem[1821] = 8'h00;
    green_mem[1822] = 8'h00;
    green_mem[1823] = 8'h00;
    green_mem[1824] = 8'h00;
    green_mem[1825] = 8'h00;
    green_mem[1826] = 8'h00;
    green_mem[1827] = 8'h00;
    green_mem[1828] = 8'h00;
    green_mem[1829] = 8'h00;
    green_mem[1830] = 8'h00;
    green_mem[1831] = 8'h00;
    green_mem[1832] = 8'h00;
    green_mem[1833] = 8'h00;
    green_mem[1834] = 8'h00;
    green_mem[1835] = 8'h00;
    green_mem[1836] = 8'h00;
    green_mem[1837] = 8'h00;
    green_mem[1838] = 8'h00;
    green_mem[1839] = 8'h00;
    green_mem[1840] = 8'h00;
    green_mem[1841] = 8'h00;
    green_mem[1842] = 8'h00;
    green_mem[1843] = 8'h00;
    green_mem[1844] = 8'h00;
    green_mem[1845] = 8'h00;
    green_mem[1846] = 8'h00;
    green_mem[1847] = 8'h00;
    green_mem[1848] = 8'h00;
    green_mem[1849] = 8'h00;
    green_mem[1850] = 8'h00;
    green_mem[1851] = 8'h00;
    green_mem[1852] = 8'h00;
    green_mem[1853] = 8'h00;
    green_mem[1854] = 8'h00;
    green_mem[1855] = 8'h00;
    green_mem[1856] = 8'h00;
    green_mem[1857] = 8'h00;
    green_mem[1858] = 8'h00;
    green_mem[1859] = 8'h00;
    green_mem[1860] = 8'h00;
    green_mem[1861] = 8'h00;
    green_mem[1862] = 8'h00;
    green_mem[1863] = 8'h00;
    green_mem[1864] = 8'h00;
    green_mem[1865] = 8'h00;
    green_mem[1866] = 8'h00;
    green_mem[1867] = 8'h00;
    green_mem[1868] = 8'h00;
    green_mem[1869] = 8'h00;
    green_mem[1870] = 8'h00;
    green_mem[1871] = 8'h00;
    green_mem[1872] = 8'h00;
    green_mem[1873] = 8'h00;
    green_mem[1874] = 8'h00;
    green_mem[1875] = 8'h00;
    green_mem[1876] = 8'h00;
    green_mem[1877] = 8'h00;
    green_mem[1878] = 8'h00;
    green_mem[1879] = 8'h00;
    green_mem[1880] = 8'h00;
    green_mem[1881] = 8'h00;
    green_mem[1882] = 8'h00;
    green_mem[1883] = 8'h00;
    green_mem[1884] = 8'h00;
    green_mem[1885] = 8'h00;
    green_mem[1886] = 8'h00;
    green_mem[1887] = 8'h00;
    green_mem[1888] = 8'h00;
    green_mem[1889] = 8'h00;
    green_mem[1890] = 8'h00;
    green_mem[1891] = 8'h00;
    green_mem[1892] = 8'h00;
    green_mem[1893] = 8'h00;
    green_mem[1894] = 8'h00;
    green_mem[1895] = 8'h00;
    green_mem[1896] = 8'h00;
    green_mem[1897] = 8'h00;
    green_mem[1898] = 8'h00;
    green_mem[1899] = 8'h00;
    green_mem[1900] = 8'h00;
    green_mem[1901] = 8'h00;
    green_mem[1902] = 8'h00;
    green_mem[1903] = 8'h00;
    green_mem[1904] = 8'h00;
    green_mem[1905] = 8'h00;
    green_mem[1906] = 8'h00;
    green_mem[1907] = 8'h00;
    green_mem[1908] = 8'h00;
    green_mem[1909] = 8'h00;
    green_mem[1910] = 8'h00;
    green_mem[1911] = 8'h00;
    green_mem[1912] = 8'h00;
    green_mem[1913] = 8'h00;
    green_mem[1914] = 8'h00;
    green_mem[1915] = 8'h00;
    green_mem[1916] = 8'h00;
    green_mem[1917] = 8'h00;
    green_mem[1918] = 8'h00;
    green_mem[1919] = 8'h00;
    green_mem[1920] = 8'h00;
    green_mem[1921] = 8'h00;
    green_mem[1922] = 8'h00;
    green_mem[1923] = 8'h00;
    green_mem[1924] = 8'h00;
    green_mem[1925] = 8'h00;
    green_mem[1926] = 8'h00;
    green_mem[1927] = 8'h00;
    green_mem[1928] = 8'h00;
    green_mem[1929] = 8'h00;
    green_mem[1930] = 8'h00;
    green_mem[1931] = 8'h00;
    green_mem[1932] = 8'h00;
    green_mem[1933] = 8'h00;
    green_mem[1934] = 8'h00;
    green_mem[1935] = 8'h00;
    green_mem[1936] = 8'h00;
    green_mem[1937] = 8'h00;
    green_mem[1938] = 8'h00;
    green_mem[1939] = 8'h00;
    green_mem[1940] = 8'h00;
    green_mem[1941] = 8'h00;
    green_mem[1942] = 8'h00;
    green_mem[1943] = 8'h00;
    green_mem[1944] = 8'h00;
    green_mem[1945] = 8'h00;
    green_mem[1946] = 8'h00;
    green_mem[1947] = 8'h00;
    green_mem[1948] = 8'h00;
    green_mem[1949] = 8'h00;
    green_mem[1950] = 8'h00;
    green_mem[1951] = 8'h00;
    green_mem[1952] = 8'h00;
    green_mem[1953] = 8'h00;
    green_mem[1954] = 8'h00;
    green_mem[1955] = 8'h00;
    green_mem[1956] = 8'h00;
    green_mem[1957] = 8'h00;
    green_mem[1958] = 8'h00;
    green_mem[1959] = 8'h00;
    green_mem[1960] = 8'h00;
    green_mem[1961] = 8'h00;
    green_mem[1962] = 8'h00;
    green_mem[1963] = 8'h00;
    green_mem[1964] = 8'h00;
    green_mem[1965] = 8'h00;
    green_mem[1966] = 8'h00;
    green_mem[1967] = 8'h00;
    green_mem[1968] = 8'h00;
    green_mem[1969] = 8'h00;
    green_mem[1970] = 8'h00;
    green_mem[1971] = 8'h00;
    green_mem[1972] = 8'h00;
    green_mem[1973] = 8'h00;
    green_mem[1974] = 8'h00;
    green_mem[1975] = 8'h00;
    green_mem[1976] = 8'h00;
    green_mem[1977] = 8'h00;
    green_mem[1978] = 8'h00;
    green_mem[1979] = 8'h00;
    green_mem[1980] = 8'h00;
    green_mem[1981] = 8'h00;
    green_mem[1982] = 8'h00;
    green_mem[1983] = 8'h00;
    green_mem[1984] = 8'h00;
    green_mem[1985] = 8'h00;
    green_mem[1986] = 8'h00;
    green_mem[1987] = 8'h00;
    green_mem[1988] = 8'h00;
    green_mem[1989] = 8'h00;
    green_mem[1990] = 8'h00;
    green_mem[1991] = 8'h00;
    green_mem[1992] = 8'h00;
    green_mem[1993] = 8'h00;
    green_mem[1994] = 8'h00;
    green_mem[1995] = 8'h00;
    green_mem[1996] = 8'h00;
    green_mem[1997] = 8'h00;
    green_mem[1998] = 8'h00;
    green_mem[1999] = 8'h00;
    green_mem[2000] = 8'h00;
    green_mem[2001] = 8'h00;
    green_mem[2002] = 8'h00;
    green_mem[2003] = 8'h00;
    green_mem[2004] = 8'h00;
    green_mem[2005] = 8'h00;
    green_mem[2006] = 8'h00;
    green_mem[2007] = 8'h00;
    green_mem[2008] = 8'h00;
    green_mem[2009] = 8'h00;
    green_mem[2010] = 8'h00;
    green_mem[2011] = 8'h00;
    green_mem[2012] = 8'h00;
    green_mem[2013] = 8'h00;
    green_mem[2014] = 8'h00;
    green_mem[2015] = 8'h00;
    green_mem[2016] = 8'h00;
    green_mem[2017] = 8'h00;
    green_mem[2018] = 8'h00;
    green_mem[2019] = 8'h00;
    green_mem[2020] = 8'h00;
    green_mem[2021] = 8'h00;
    green_mem[2022] = 8'h00;
    green_mem[2023] = 8'h00;
    green_mem[2024] = 8'h00;
    green_mem[2025] = 8'h00;
    green_mem[2026] = 8'h00;
    green_mem[2027] = 8'h00;
    green_mem[2028] = 8'h00;
    green_mem[2029] = 8'h00;
    green_mem[2030] = 8'h00;
    green_mem[2031] = 8'h00;
    green_mem[2032] = 8'h00;
    green_mem[2033] = 8'h00;
    green_mem[2034] = 8'h00;
    green_mem[2035] = 8'h00;
    green_mem[2036] = 8'h00;
    green_mem[2037] = 8'h00;
    green_mem[2038] = 8'h00;
    green_mem[2039] = 8'h00;
    green_mem[2040] = 8'h00;
    green_mem[2041] = 8'h00;
    green_mem[2042] = 8'h00;
    green_mem[2043] = 8'h00;
    green_mem[2044] = 8'h00;
    green_mem[2045] = 8'h00;
    green_mem[2046] = 8'h00;
    green_mem[2047] = 8'h00;
    blue_mem[0] = 8'h00;
    blue_mem[1] = 8'h00;
    blue_mem[2] = 8'h00;
    blue_mem[3] = 8'h00;
    blue_mem[4] = 8'h00;
    blue_mem[5] = 8'h00;
    blue_mem[6] = 8'h00;
    blue_mem[7] = 8'h00;
    blue_mem[8] = 8'h00;
    blue_mem[9] = 8'h00;
    blue_mem[10] = 8'h00;
    blue_mem[11] = 8'h00;
    blue_mem[12] = 8'h00;
    blue_mem[13] = 8'h00;
    blue_mem[14] = 8'h00;
    blue_mem[15] = 8'h00;
    blue_mem[16] = 8'h00;
    blue_mem[17] = 8'h00;
    blue_mem[18] = 8'h00;
    blue_mem[19] = 8'h00;
    blue_mem[20] = 8'h00;
    blue_mem[21] = 8'h00;
    blue_mem[22] = 8'h00;
    blue_mem[23] = 8'h00;
    blue_mem[24] = 8'h00;
    blue_mem[25] = 8'h00;
    blue_mem[26] = 8'h00;
    blue_mem[27] = 8'h00;
    blue_mem[28] = 8'h00;
    blue_mem[29] = 8'h00;
    blue_mem[30] = 8'h00;
    blue_mem[31] = 8'h00;
    blue_mem[32] = 8'h00;
    blue_mem[33] = 8'h00;
    blue_mem[34] = 8'h00;
    blue_mem[35] = 8'h00;
    blue_mem[36] = 8'h00;
    blue_mem[37] = 8'h00;
    blue_mem[38] = 8'h00;
    blue_mem[39] = 8'h00;
    blue_mem[40] = 8'h00;
    blue_mem[41] = 8'h00;
    blue_mem[42] = 8'h00;
    blue_mem[43] = 8'h00;
    blue_mem[44] = 8'h00;
    blue_mem[45] = 8'h00;
    blue_mem[46] = 8'h00;
    blue_mem[47] = 8'h00;
    blue_mem[48] = 8'h00;
    blue_mem[49] = 8'h00;
    blue_mem[50] = 8'h00;
    blue_mem[51] = 8'h00;
    blue_mem[52] = 8'h00;
    blue_mem[53] = 8'h00;
    blue_mem[54] = 8'h00;
    blue_mem[55] = 8'h00;
    blue_mem[56] = 8'h00;
    blue_mem[57] = 8'h00;
    blue_mem[58] = 8'h00;
    blue_mem[59] = 8'h00;
    blue_mem[60] = 8'h00;
    blue_mem[61] = 8'h00;
    blue_mem[62] = 8'h00;
    blue_mem[63] = 8'h00;
    blue_mem[64] = 8'h00;
    blue_mem[65] = 8'h00;
    blue_mem[66] = 8'h00;
    blue_mem[67] = 8'h00;
    blue_mem[68] = 8'h00;
    blue_mem[69] = 8'h00;
    blue_mem[70] = 8'h00;
    blue_mem[71] = 8'h00;
    blue_mem[72] = 8'h00;
    blue_mem[73] = 8'h00;
    blue_mem[74] = 8'h00;
    blue_mem[75] = 8'h00;
    blue_mem[76] = 8'h00;
    blue_mem[77] = 8'h00;
    blue_mem[78] = 8'h00;
    blue_mem[79] = 8'h00;
    blue_mem[80] = 8'h00;
    blue_mem[81] = 8'h00;
    blue_mem[82] = 8'h00;
    blue_mem[83] = 8'h00;
    blue_mem[84] = 8'h00;
    blue_mem[85] = 8'h00;
    blue_mem[86] = 8'h00;
    blue_mem[87] = 8'h00;
    blue_mem[88] = 8'h00;
    blue_mem[89] = 8'h00;
    blue_mem[90] = 8'h00;
    blue_mem[91] = 8'h00;
    blue_mem[92] = 8'h00;
    blue_mem[93] = 8'h00;
    blue_mem[94] = 8'h00;
    blue_mem[95] = 8'h00;
    blue_mem[96] = 8'h00;
    blue_mem[97] = 8'h00;
    blue_mem[98] = 8'h00;
    blue_mem[99] = 8'h00;
    blue_mem[100] = 8'h00;
    blue_mem[101] = 8'h00;
    blue_mem[102] = 8'h00;
    blue_mem[103] = 8'h00;
    blue_mem[104] = 8'h00;
    blue_mem[105] = 8'h00;
    blue_mem[106] = 8'h00;
    blue_mem[107] = 8'h00;
    blue_mem[108] = 8'h00;
    blue_mem[109] = 8'h00;
    blue_mem[110] = 8'h00;
    blue_mem[111] = 8'h00;
    blue_mem[112] = 8'h00;
    blue_mem[113] = 8'h00;
    blue_mem[114] = 8'h00;
    blue_mem[115] = 8'h00;
    blue_mem[116] = 8'h00;
    blue_mem[117] = 8'h00;
    blue_mem[118] = 8'h00;
    blue_mem[119] = 8'h00;
    blue_mem[120] = 8'h00;
    blue_mem[121] = 8'h00;
    blue_mem[122] = 8'h00;
    blue_mem[123] = 8'h00;
    blue_mem[124] = 8'h00;
    blue_mem[125] = 8'h00;
    blue_mem[126] = 8'h00;
    blue_mem[127] = 8'h00;
    blue_mem[128] = 8'h00;
    blue_mem[129] = 8'h00;
    blue_mem[130] = 8'h00;
    blue_mem[131] = 8'h00;
    blue_mem[132] = 8'h00;
    blue_mem[133] = 8'h00;
    blue_mem[134] = 8'h00;
    blue_mem[135] = 8'h00;
    blue_mem[136] = 8'h00;
    blue_mem[137] = 8'h00;
    blue_mem[138] = 8'h00;
    blue_mem[139] = 8'h00;
    blue_mem[140] = 8'h00;
    blue_mem[141] = 8'h00;
    blue_mem[142] = 8'h00;
    blue_mem[143] = 8'h00;
    blue_mem[144] = 8'h00;
    blue_mem[145] = 8'h00;
    blue_mem[146] = 8'h00;
    blue_mem[147] = 8'h00;
    blue_mem[148] = 8'h00;
    blue_mem[149] = 8'h00;
    blue_mem[150] = 8'h00;
    blue_mem[151] = 8'h00;
    blue_mem[152] = 8'h00;
    blue_mem[153] = 8'h00;
    blue_mem[154] = 8'h00;
    blue_mem[155] = 8'h00;
    blue_mem[156] = 8'h00;
    blue_mem[157] = 8'h00;
    blue_mem[158] = 8'h00;
    blue_mem[159] = 8'h00;
    blue_mem[160] = 8'h00;
    blue_mem[161] = 8'h00;
    blue_mem[162] = 8'h00;
    blue_mem[163] = 8'h00;
    blue_mem[164] = 8'h00;
    blue_mem[165] = 8'h00;
    blue_mem[166] = 8'h00;
    blue_mem[167] = 8'h00;
    blue_mem[168] = 8'h00;
    blue_mem[169] = 8'h00;
    blue_mem[170] = 8'h00;
    blue_mem[171] = 8'h00;
    blue_mem[172] = 8'h00;
    blue_mem[173] = 8'h00;
    blue_mem[174] = 8'h00;
    blue_mem[175] = 8'h00;
    blue_mem[176] = 8'h00;
    blue_mem[177] = 8'h00;
    blue_mem[178] = 8'h00;
    blue_mem[179] = 8'h00;
    blue_mem[180] = 8'h00;
    blue_mem[181] = 8'h00;
    blue_mem[182] = 8'h00;
    blue_mem[183] = 8'h00;
    blue_mem[184] = 8'h00;
    blue_mem[185] = 8'h00;
    blue_mem[186] = 8'h00;
    blue_mem[187] = 8'h00;
    blue_mem[188] = 8'h00;
    blue_mem[189] = 8'h00;
    blue_mem[190] = 8'h00;
    blue_mem[191] = 8'h00;
    blue_mem[192] = 8'h00;
    blue_mem[193] = 8'h00;
    blue_mem[194] = 8'h00;
    blue_mem[195] = 8'h00;
    blue_mem[196] = 8'h00;
    blue_mem[197] = 8'h00;
    blue_mem[198] = 8'h00;
    blue_mem[199] = 8'h00;
    blue_mem[200] = 8'h00;
    blue_mem[201] = 8'h00;
    blue_mem[202] = 8'h00;
    blue_mem[203] = 8'h00;
    blue_mem[204] = 8'h00;
    blue_mem[205] = 8'h00;
    blue_mem[206] = 8'h00;
    blue_mem[207] = 8'h00;
    blue_mem[208] = 8'h00;
    blue_mem[209] = 8'h00;
    blue_mem[210] = 8'h00;
    blue_mem[211] = 8'h00;
    blue_mem[212] = 8'h00;
    blue_mem[213] = 8'h00;
    blue_mem[214] = 8'h00;
    blue_mem[215] = 8'h00;
    blue_mem[216] = 8'h00;
    blue_mem[217] = 8'h00;
    blue_mem[218] = 8'h00;
    blue_mem[219] = 8'h00;
    blue_mem[220] = 8'h00;
    blue_mem[221] = 8'h00;
    blue_mem[222] = 8'h00;
    blue_mem[223] = 8'h00;
    blue_mem[224] = 8'h00;
    blue_mem[225] = 8'h00;
    blue_mem[226] = 8'h00;
    blue_mem[227] = 8'h00;
    blue_mem[228] = 8'h00;
    blue_mem[229] = 8'h00;
    blue_mem[230] = 8'h00;
    blue_mem[231] = 8'h00;
    blue_mem[232] = 8'h00;
    blue_mem[233] = 8'h00;
    blue_mem[234] = 8'h00;
    blue_mem[235] = 8'h00;
    blue_mem[236] = 8'h00;
    blue_mem[237] = 8'h00;
    blue_mem[238] = 8'h00;
    blue_mem[239] = 8'h00;
    blue_mem[240] = 8'h00;
    blue_mem[241] = 8'h00;
    blue_mem[242] = 8'h00;
    blue_mem[243] = 8'h00;
    blue_mem[244] = 8'h00;
    blue_mem[245] = 8'h00;
    blue_mem[246] = 8'h00;
    blue_mem[247] = 8'h00;
    blue_mem[248] = 8'h00;
    blue_mem[249] = 8'h00;
    blue_mem[250] = 8'h00;
    blue_mem[251] = 8'h00;
    blue_mem[252] = 8'h00;
    blue_mem[253] = 8'h00;
    blue_mem[254] = 8'h00;
    blue_mem[255] = 8'h00;
    blue_mem[256] = 8'h00;
    blue_mem[257] = 8'h00;
    blue_mem[258] = 8'h00;
    blue_mem[259] = 8'h00;
    blue_mem[260] = 8'h00;
    blue_mem[261] = 8'h00;
    blue_mem[262] = 8'h00;
    blue_mem[263] = 8'h00;
    blue_mem[264] = 8'h10;
    blue_mem[265] = 8'h00;
    blue_mem[266] = 8'h00;
    blue_mem[267] = 8'h00;
    blue_mem[268] = 8'h00;
    blue_mem[269] = 8'h00;
    blue_mem[270] = 8'h00;
    blue_mem[271] = 8'h00;
    blue_mem[272] = 8'h00;
    blue_mem[273] = 8'h00;
    blue_mem[274] = 8'h00;
    blue_mem[275] = 8'h00;
    blue_mem[276] = 8'h00;
    blue_mem[277] = 8'h00;
    blue_mem[278] = 8'h00;
    blue_mem[279] = 8'hd8;
    blue_mem[280] = 8'hfd;
    blue_mem[281] = 8'h03;
    blue_mem[282] = 8'h00;
    blue_mem[283] = 8'h00;
    blue_mem[284] = 8'h00;
    blue_mem[285] = 8'h00;
    blue_mem[286] = 8'h00;
    blue_mem[287] = 8'h00;
    blue_mem[288] = 8'h00;
    blue_mem[289] = 8'h00;
    blue_mem[290] = 8'h00;
    blue_mem[291] = 8'h00;
    blue_mem[292] = 8'h00;
    blue_mem[293] = 8'h00;
    blue_mem[294] = 8'hb8;
    blue_mem[295] = 8'hff;
    blue_mem[296] = 8'hff;
    blue_mem[297] = 8'h3b;
    blue_mem[298] = 8'h00;
    blue_mem[299] = 8'h00;
    blue_mem[300] = 8'h00;
    blue_mem[301] = 8'h00;
    blue_mem[302] = 8'h00;
    blue_mem[303] = 8'h00;
    blue_mem[304] = 8'h00;
    blue_mem[305] = 8'h00;
    blue_mem[306] = 8'h00;
    blue_mem[307] = 8'h00;
    blue_mem[308] = 8'h00;
    blue_mem[309] = 8'h00;
    blue_mem[310] = 8'hfc;
    blue_mem[311] = 8'hff;
    blue_mem[312] = 8'hff;
    blue_mem[313] = 8'hfb;
    blue_mem[314] = 8'h03;
    blue_mem[315] = 8'h00;
    blue_mem[316] = 8'h00;
    blue_mem[317] = 8'h00;
    blue_mem[318] = 8'h00;
    blue_mem[319] = 8'h00;
    blue_mem[320] = 8'h00;
    blue_mem[321] = 8'h00;
    blue_mem[322] = 8'h00;
    blue_mem[323] = 8'h00;
    blue_mem[324] = 8'h00;
    blue_mem[325] = 8'hc0;
    blue_mem[326] = 8'hff;
    blue_mem[327] = 8'hff;
    blue_mem[328] = 8'hff;
    blue_mem[329] = 8'hff;
    blue_mem[330] = 8'h03;
    blue_mem[331] = 8'h00;
    blue_mem[332] = 8'h00;
    blue_mem[333] = 8'h00;
    blue_mem[334] = 8'h00;
    blue_mem[335] = 8'h00;
    blue_mem[336] = 8'h00;
    blue_mem[337] = 8'h00;
    blue_mem[338] = 8'h00;
    blue_mem[339] = 8'h00;
    blue_mem[340] = 8'h00;
    blue_mem[341] = 8'he0;
    blue_mem[342] = 8'hff;
    blue_mem[343] = 8'hff;
    blue_mem[344] = 8'hff;
    blue_mem[345] = 8'hff;
    blue_mem[346] = 8'h17;
    blue_mem[347] = 8'h00;
    blue_mem[348] = 8'h00;
    blue_mem[349] = 8'h00;
    blue_mem[350] = 8'h00;
    blue_mem[351] = 8'h00;
    blue_mem[352] = 8'h00;
    blue_mem[353] = 8'h00;
    blue_mem[354] = 8'h00;
    blue_mem[355] = 8'h00;
    blue_mem[356] = 8'h00;
    blue_mem[357] = 8'hfc;
    blue_mem[358] = 8'hff;
    blue_mem[359] = 8'hff;
    blue_mem[360] = 8'hff;
    blue_mem[361] = 8'hff;
    blue_mem[362] = 8'h3f;
    blue_mem[363] = 8'h00;
    blue_mem[364] = 8'h00;
    blue_mem[365] = 8'h00;
    blue_mem[366] = 8'h00;
    blue_mem[367] = 8'h00;
    blue_mem[368] = 8'h00;
    blue_mem[369] = 8'h00;
    blue_mem[370] = 8'h00;
    blue_mem[371] = 8'h00;
    blue_mem[372] = 8'h00;
    blue_mem[373] = 8'hfc;
    blue_mem[374] = 8'hff;
    blue_mem[375] = 8'hff;
    blue_mem[376] = 8'hff;
    blue_mem[377] = 8'hff;
    blue_mem[378] = 8'h3f;
    blue_mem[379] = 8'h00;
    blue_mem[380] = 8'h00;
    blue_mem[381] = 8'h00;
    blue_mem[382] = 8'h00;
    blue_mem[383] = 8'h00;
    blue_mem[384] = 8'h00;
    blue_mem[385] = 8'h00;
    blue_mem[386] = 8'h00;
    blue_mem[387] = 8'h00;
    blue_mem[388] = 8'hc0;
    blue_mem[389] = 8'hff;
    blue_mem[390] = 8'hff;
    blue_mem[391] = 8'hff;
    blue_mem[392] = 8'hff;
    blue_mem[393] = 8'hff;
    blue_mem[394] = 8'hff;
    blue_mem[395] = 8'h07;
    blue_mem[396] = 8'h00;
    blue_mem[397] = 8'h00;
    blue_mem[398] = 8'h00;
    blue_mem[399] = 8'h00;
    blue_mem[400] = 8'h00;
    blue_mem[401] = 8'h00;
    blue_mem[402] = 8'h00;
    blue_mem[403] = 8'h00;
    blue_mem[404] = 8'hc0;
    blue_mem[405] = 8'hff;
    blue_mem[406] = 8'hff;
    blue_mem[407] = 8'hff;
    blue_mem[408] = 8'hff;
    blue_mem[409] = 8'hff;
    blue_mem[410] = 8'hff;
    blue_mem[411] = 8'h0f;
    blue_mem[412] = 8'h00;
    blue_mem[413] = 8'h00;
    blue_mem[414] = 8'h00;
    blue_mem[415] = 8'h00;
    blue_mem[416] = 8'h00;
    blue_mem[417] = 8'h00;
    blue_mem[418] = 8'h00;
    blue_mem[419] = 8'h00;
    blue_mem[420] = 8'hf8;
    blue_mem[421] = 8'hff;
    blue_mem[422] = 8'hff;
    blue_mem[423] = 8'hff;
    blue_mem[424] = 8'hff;
    blue_mem[425] = 8'hff;
    blue_mem[426] = 8'hff;
    blue_mem[427] = 8'h0f;
    blue_mem[428] = 8'h00;
    blue_mem[429] = 8'h00;
    blue_mem[430] = 8'h00;
    blue_mem[431] = 8'h00;
    blue_mem[432] = 8'h00;
    blue_mem[433] = 8'h00;
    blue_mem[434] = 8'h00;
    blue_mem[435] = 8'h00;
    blue_mem[436] = 8'hf8;
    blue_mem[437] = 8'hff;
    blue_mem[438] = 8'hbf;
    blue_mem[439] = 8'hff;
    blue_mem[440] = 8'hff;
    blue_mem[441] = 8'hff;
    blue_mem[442] = 8'hff;
    blue_mem[443] = 8'h3f;
    blue_mem[444] = 8'h00;
    blue_mem[445] = 8'h00;
    blue_mem[446] = 8'h00;
    blue_mem[447] = 8'h00;
    blue_mem[448] = 8'h00;
    blue_mem[449] = 8'h00;
    blue_mem[450] = 8'h00;
    blue_mem[451] = 8'h00;
    blue_mem[452] = 8'hf8;
    blue_mem[453] = 8'hff;
    blue_mem[454] = 8'hff;
    blue_mem[455] = 8'hff;
    blue_mem[456] = 8'hff;
    blue_mem[457] = 8'hff;
    blue_mem[458] = 8'hff;
    blue_mem[459] = 8'h7f;
    blue_mem[460] = 8'h00;
    blue_mem[461] = 8'h00;
    blue_mem[462] = 8'h00;
    blue_mem[463] = 8'h00;
    blue_mem[464] = 8'h00;
    blue_mem[465] = 8'h00;
    blue_mem[466] = 8'h00;
    blue_mem[467] = 8'h00;
    blue_mem[468] = 8'hfe;
    blue_mem[469] = 8'hff;
    blue_mem[470] = 8'hff;
    blue_mem[471] = 8'hff;
    blue_mem[472] = 8'hff;
    blue_mem[473] = 8'hff;
    blue_mem[474] = 8'hff;
    blue_mem[475] = 8'hff;
    blue_mem[476] = 8'h01;
    blue_mem[477] = 8'h00;
    blue_mem[478] = 8'h00;
    blue_mem[479] = 8'h00;
    blue_mem[480] = 8'h00;
    blue_mem[481] = 8'h00;
    blue_mem[482] = 8'h00;
    blue_mem[483] = 8'h80;
    blue_mem[484] = 8'hff;
    blue_mem[485] = 8'hfe;
    blue_mem[486] = 8'hff;
    blue_mem[487] = 8'hff;
    blue_mem[488] = 8'hff;
    blue_mem[489] = 8'hff;
    blue_mem[490] = 8'hff;
    blue_mem[491] = 8'hff;
    blue_mem[492] = 8'h01;
    blue_mem[493] = 8'h00;
    blue_mem[494] = 8'h00;
    blue_mem[495] = 8'h00;
    blue_mem[496] = 8'h00;
    blue_mem[497] = 8'h00;
    blue_mem[498] = 8'h00;
    blue_mem[499] = 8'hc0;
    blue_mem[500] = 8'hff;
    blue_mem[501] = 8'hff;
    blue_mem[502] = 8'hff;
    blue_mem[503] = 8'hff;
    blue_mem[504] = 8'hff;
    blue_mem[505] = 8'hff;
    blue_mem[506] = 8'hff;
    blue_mem[507] = 8'hff;
    blue_mem[508] = 8'h03;
    blue_mem[509] = 8'h00;
    blue_mem[510] = 8'h00;
    blue_mem[511] = 8'h00;
    blue_mem[512] = 8'h00;
    blue_mem[513] = 8'h00;
    blue_mem[514] = 8'h00;
    blue_mem[515] = 8'hc0;
    blue_mem[516] = 8'hff;
    blue_mem[517] = 8'hff;
    blue_mem[518] = 8'hff;
    blue_mem[519] = 8'hff;
    blue_mem[520] = 8'hff;
    blue_mem[521] = 8'hff;
    blue_mem[522] = 8'hff;
    blue_mem[523] = 8'hff;
    blue_mem[524] = 8'h07;
    blue_mem[525] = 8'h00;
    blue_mem[526] = 8'h00;
    blue_mem[527] = 8'h00;
    blue_mem[528] = 8'h00;
    blue_mem[529] = 8'h00;
    blue_mem[530] = 8'h00;
    blue_mem[531] = 8'hc0;
    blue_mem[532] = 8'hff;
    blue_mem[533] = 8'hf7;
    blue_mem[534] = 8'hff;
    blue_mem[535] = 8'hff;
    blue_mem[536] = 8'hff;
    blue_mem[537] = 8'hff;
    blue_mem[538] = 8'hff;
    blue_mem[539] = 8'hff;
    blue_mem[540] = 8'h0f;
    blue_mem[541] = 8'h00;
    blue_mem[542] = 8'h00;
    blue_mem[543] = 8'h00;
    blue_mem[544] = 8'h00;
    blue_mem[545] = 8'h00;
    blue_mem[546] = 8'h00;
    blue_mem[547] = 8'hf8;
    blue_mem[548] = 8'hff;
    blue_mem[549] = 8'hff;
    blue_mem[550] = 8'hdf;
    blue_mem[551] = 8'hff;
    blue_mem[552] = 8'hff;
    blue_mem[553] = 8'hff;
    blue_mem[554] = 8'hff;
    blue_mem[555] = 8'hff;
    blue_mem[556] = 8'h1f;
    blue_mem[557] = 8'h00;
    blue_mem[558] = 8'h00;
    blue_mem[559] = 8'h00;
    blue_mem[560] = 8'h00;
    blue_mem[561] = 8'h00;
    blue_mem[562] = 8'h00;
    blue_mem[563] = 8'hf8;
    blue_mem[564] = 8'hff;
    blue_mem[565] = 8'hff;
    blue_mem[566] = 8'hfd;
    blue_mem[567] = 8'hff;
    blue_mem[568] = 8'hff;
    blue_mem[569] = 8'hff;
    blue_mem[570] = 8'hff;
    blue_mem[571] = 8'hfe;
    blue_mem[572] = 8'h1d;
    blue_mem[573] = 8'h00;
    blue_mem[574] = 8'h00;
    blue_mem[575] = 8'h00;
    blue_mem[576] = 8'h00;
    blue_mem[577] = 8'h00;
    blue_mem[578] = 8'h00;
    blue_mem[579] = 8'hf0;
    blue_mem[580] = 8'hff;
    blue_mem[581] = 8'hff;
    blue_mem[582] = 8'hff;
    blue_mem[583] = 8'hff;
    blue_mem[584] = 8'hff;
    blue_mem[585] = 8'hff;
    blue_mem[586] = 8'hff;
    blue_mem[587] = 8'hff;
    blue_mem[588] = 8'h7b;
    blue_mem[589] = 8'h00;
    blue_mem[590] = 8'h00;
    blue_mem[591] = 8'h00;
    blue_mem[592] = 8'h00;
    blue_mem[593] = 8'h00;
    blue_mem[594] = 8'h00;
    blue_mem[595] = 8'hfe;
    blue_mem[596] = 8'hbf;
    blue_mem[597] = 8'hff;
    blue_mem[598] = 8'h1f;
    blue_mem[599] = 8'hff;
    blue_mem[600] = 8'hff;
    blue_mem[601] = 8'h0f;
    blue_mem[602] = 8'hc0;
    blue_mem[603] = 8'hff;
    blue_mem[604] = 8'hff;
    blue_mem[605] = 8'h00;
    blue_mem[606] = 8'h00;
    blue_mem[607] = 8'h00;
    blue_mem[608] = 8'h00;
    blue_mem[609] = 8'h00;
    blue_mem[610] = 8'h00;
    blue_mem[611] = 8'hfe;
    blue_mem[612] = 8'hfd;
    blue_mem[613] = 8'hff;
    blue_mem[614] = 8'h07;
    blue_mem[615] = 8'hff;
    blue_mem[616] = 8'hff;
    blue_mem[617] = 8'h00;
    blue_mem[618] = 8'h00;
    blue_mem[619] = 8'hfc;
    blue_mem[620] = 8'hff;
    blue_mem[621] = 8'h00;
    blue_mem[622] = 8'h00;
    blue_mem[623] = 8'h00;
    blue_mem[624] = 8'h00;
    blue_mem[625] = 8'h00;
    blue_mem[626] = 8'h00;
    blue_mem[627] = 8'hfe;
    blue_mem[628] = 8'hff;
    blue_mem[629] = 8'hff;
    blue_mem[630] = 8'h03;
    blue_mem[631] = 8'hff;
    blue_mem[632] = 8'hff;
    blue_mem[633] = 8'h00;
    blue_mem[634] = 8'h00;
    blue_mem[635] = 8'hf0;
    blue_mem[636] = 8'hff;
    blue_mem[637] = 8'h00;
    blue_mem[638] = 8'h00;
    blue_mem[639] = 8'h00;
    blue_mem[640] = 8'h00;
    blue_mem[641] = 8'h00;
    blue_mem[642] = 8'h80;
    blue_mem[643] = 8'hff;
    blue_mem[644] = 8'hff;
    blue_mem[645] = 8'hff;
    blue_mem[646] = 8'h80;
    blue_mem[647] = 8'hff;
    blue_mem[648] = 8'h1f;
    blue_mem[649] = 8'h00;
    blue_mem[650] = 8'h00;
    blue_mem[651] = 8'hf0;
    blue_mem[652] = 8'hff;
    blue_mem[653] = 8'h01;
    blue_mem[654] = 8'h00;
    blue_mem[655] = 8'h00;
    blue_mem[656] = 8'h00;
    blue_mem[657] = 8'h00;
    blue_mem[658] = 8'h80;
    blue_mem[659] = 8'hff;
    blue_mem[660] = 8'hef;
    blue_mem[661] = 8'hff;
    blue_mem[662] = 8'h00;
    blue_mem[663] = 8'hff;
    blue_mem[664] = 8'h1b;
    blue_mem[665] = 8'hf0;
    blue_mem[666] = 8'h00;
    blue_mem[667] = 8'he0;
    blue_mem[668] = 8'hff;
    blue_mem[669] = 8'h01;
    blue_mem[670] = 8'h00;
    blue_mem[671] = 8'h00;
    blue_mem[672] = 8'h00;
    blue_mem[673] = 8'h00;
    blue_mem[674] = 8'hc0;
    blue_mem[675] = 8'hff;
    blue_mem[676] = 8'hef;
    blue_mem[677] = 8'hfe;
    blue_mem[678] = 8'h00;
    blue_mem[679] = 8'hff;
    blue_mem[680] = 8'h03;
    blue_mem[681] = 8'hf8;
    blue_mem[682] = 8'h07;
    blue_mem[683] = 8'he0;
    blue_mem[684] = 8'hff;
    blue_mem[685] = 8'h03;
    blue_mem[686] = 8'h00;
    blue_mem[687] = 8'h00;
    blue_mem[688] = 8'h00;
    blue_mem[689] = 8'h00;
    blue_mem[690] = 8'hc0;
    blue_mem[691] = 8'hbf;
    blue_mem[692] = 8'hff;
    blue_mem[693] = 8'h3f;
    blue_mem[694] = 8'h80;
    blue_mem[695] = 8'hef;
    blue_mem[696] = 8'h07;
    blue_mem[697] = 8'hfc;
    blue_mem[698] = 8'h3f;
    blue_mem[699] = 8'he0;
    blue_mem[700] = 8'hff;
    blue_mem[701] = 8'h07;
    blue_mem[702] = 8'h00;
    blue_mem[703] = 8'h00;
    blue_mem[704] = 8'h00;
    blue_mem[705] = 8'h00;
    blue_mem[706] = 8'he0;
    blue_mem[707] = 8'hff;
    blue_mem[708] = 8'hff;
    blue_mem[709] = 8'h3f;
    blue_mem[710] = 8'h80;
    blue_mem[711] = 8'hff;
    blue_mem[712] = 8'h03;
    blue_mem[713] = 8'hfe;
    blue_mem[714] = 8'h7f;
    blue_mem[715] = 8'h80;
    blue_mem[716] = 8'hff;
    blue_mem[717] = 8'h07;
    blue_mem[718] = 8'h00;
    blue_mem[719] = 8'h00;
    blue_mem[720] = 8'h00;
    blue_mem[721] = 8'h00;
    blue_mem[722] = 8'hc0;
    blue_mem[723] = 8'hff;
    blue_mem[724] = 8'hff;
    blue_mem[725] = 8'h0f;
    blue_mem[726] = 8'h80;
    blue_mem[727] = 8'hff;
    blue_mem[728] = 8'h03;
    blue_mem[729] = 8'hff;
    blue_mem[730] = 8'h7f;
    blue_mem[731] = 8'h00;
    blue_mem[732] = 8'hff;
    blue_mem[733] = 8'h0f;
    blue_mem[734] = 8'h00;
    blue_mem[735] = 8'h00;
    blue_mem[736] = 8'h00;
    blue_mem[737] = 8'h00;
    blue_mem[738] = 8'hf0;
    blue_mem[739] = 8'hfd;
    blue_mem[740] = 8'hdf;
    blue_mem[741] = 8'h0f;
    blue_mem[742] = 8'h80;
    blue_mem[743] = 8'hff;
    blue_mem[744] = 8'h01;
    blue_mem[745] = 8'hff;
    blue_mem[746] = 8'hff;
    blue_mem[747] = 8'h80;
    blue_mem[748] = 8'hff;
    blue_mem[749] = 8'h0f;
    blue_mem[750] = 8'h00;
    blue_mem[751] = 8'h00;
    blue_mem[752] = 8'h00;
    blue_mem[753] = 8'h00;
    blue_mem[754] = 8'hf0;
    blue_mem[755] = 8'hff;
    blue_mem[756] = 8'hff;
    blue_mem[757] = 8'h0f;
    blue_mem[758] = 8'h80;
    blue_mem[759] = 8'hff;
    blue_mem[760] = 8'h03;
    blue_mem[761] = 8'hff;
    blue_mem[762] = 8'hff;
    blue_mem[763] = 8'h00;
    blue_mem[764] = 8'hff;
    blue_mem[765] = 8'h1f;
    blue_mem[766] = 8'h00;
    blue_mem[767] = 8'h00;
    blue_mem[768] = 8'h00;
    blue_mem[769] = 8'h00;
    blue_mem[770] = 8'hf0;
    blue_mem[771] = 8'hff;
    blue_mem[772] = 8'hff;
    blue_mem[773] = 8'h01;
    blue_mem[774] = 8'hc0;
    blue_mem[775] = 8'hff;
    blue_mem[776] = 8'h01;
    blue_mem[777] = 8'hff;
    blue_mem[778] = 8'h7f;
    blue_mem[779] = 8'h00;
    blue_mem[780] = 8'hff;
    blue_mem[781] = 8'h1f;
    blue_mem[782] = 8'h00;
    blue_mem[783] = 8'h00;
    blue_mem[784] = 8'h00;
    blue_mem[785] = 8'h00;
    blue_mem[786] = 8'hf0;
    blue_mem[787] = 8'hff;
    blue_mem[788] = 8'hff;
    blue_mem[789] = 8'h61;
    blue_mem[790] = 8'hc0;
    blue_mem[791] = 8'hff;
    blue_mem[792] = 8'h01;
    blue_mem[793] = 8'hfe;
    blue_mem[794] = 8'h6f;
    blue_mem[795] = 8'h00;
    blue_mem[796] = 8'hff;
    blue_mem[797] = 8'h1f;
    blue_mem[798] = 8'h00;
    blue_mem[799] = 8'h00;
    blue_mem[800] = 8'h00;
    blue_mem[801] = 8'h00;
    blue_mem[802] = 8'hf8;
    blue_mem[803] = 8'hff;
    blue_mem[804] = 8'h3f;
    blue_mem[805] = 8'h60;
    blue_mem[806] = 8'hc0;
    blue_mem[807] = 8'hff;
    blue_mem[808] = 8'h00;
    blue_mem[809] = 8'hf8;
    blue_mem[810] = 8'hff;
    blue_mem[811] = 8'h00;
    blue_mem[812] = 8'h9f;
    blue_mem[813] = 8'h3f;
    blue_mem[814] = 8'h00;
    blue_mem[815] = 8'h00;
    blue_mem[816] = 8'h00;
    blue_mem[817] = 8'h00;
    blue_mem[818] = 8'hfc;
    blue_mem[819] = 8'hff;
    blue_mem[820] = 8'h3f;
    blue_mem[821] = 8'h70;
    blue_mem[822] = 8'he0;
    blue_mem[823] = 8'hff;
    blue_mem[824] = 8'h00;
    blue_mem[825] = 8'hb8;
    blue_mem[826] = 8'h3f;
    blue_mem[827] = 8'h00;
    blue_mem[828] = 8'hff;
    blue_mem[829] = 8'h3f;
    blue_mem[830] = 8'h00;
    blue_mem[831] = 8'h00;
    blue_mem[832] = 8'h00;
    blue_mem[833] = 8'h00;
    blue_mem[834] = 8'hfc;
    blue_mem[835] = 8'hff;
    blue_mem[836] = 8'h3f;
    blue_mem[837] = 8'h38;
    blue_mem[838] = 8'he0;
    blue_mem[839] = 8'hfe;
    blue_mem[840] = 8'h00;
    blue_mem[841] = 8'hf0;
    blue_mem[842] = 8'h3f;
    blue_mem[843] = 8'h00;
    blue_mem[844] = 8'hff;
    blue_mem[845] = 8'h3f;
    blue_mem[846] = 8'h00;
    blue_mem[847] = 8'h00;
    blue_mem[848] = 8'h00;
    blue_mem[849] = 8'h00;
    blue_mem[850] = 8'hfc;
    blue_mem[851] = 8'hff;
    blue_mem[852] = 8'h3f;
    blue_mem[853] = 8'h3c;
    blue_mem[854] = 8'he0;
    blue_mem[855] = 8'hff;
    blue_mem[856] = 8'h00;
    blue_mem[857] = 8'hf8;
    blue_mem[858] = 8'h3f;
    blue_mem[859] = 8'h80;
    blue_mem[860] = 8'hff;
    blue_mem[861] = 8'h3f;
    blue_mem[862] = 8'h00;
    blue_mem[863] = 8'h00;
    blue_mem[864] = 8'h00;
    blue_mem[865] = 8'h00;
    blue_mem[866] = 8'hf8;
    blue_mem[867] = 8'hff;
    blue_mem[868] = 8'h3f;
    blue_mem[869] = 8'h3e;
    blue_mem[870] = 8'he0;
    blue_mem[871] = 8'hff;
    blue_mem[872] = 8'h00;
    blue_mem[873] = 8'hf8;
    blue_mem[874] = 8'h3f;
    blue_mem[875] = 8'h80;
    blue_mem[876] = 8'hff;
    blue_mem[877] = 8'h3f;
    blue_mem[878] = 8'h00;
    blue_mem[879] = 8'h00;
    blue_mem[880] = 8'h00;
    blue_mem[881] = 8'h00;
    blue_mem[882] = 8'hfc;
    blue_mem[883] = 8'hff;
    blue_mem[884] = 8'hbb;
    blue_mem[885] = 8'h1f;
    blue_mem[886] = 8'hf0;
    blue_mem[887] = 8'hff;
    blue_mem[888] = 8'h00;
    blue_mem[889] = 8'hf8;
    blue_mem[890] = 8'h1d;
    blue_mem[891] = 8'h80;
    blue_mem[892] = 8'hff;
    blue_mem[893] = 8'h7f;
    blue_mem[894] = 8'h00;
    blue_mem[895] = 8'h00;
    blue_mem[896] = 8'h00;
    blue_mem[897] = 8'h00;
    blue_mem[898] = 8'hfc;
    blue_mem[899] = 8'hff;
    blue_mem[900] = 8'hff;
    blue_mem[901] = 8'h1f;
    blue_mem[902] = 8'he0;
    blue_mem[903] = 8'hff;
    blue_mem[904] = 8'h03;
    blue_mem[905] = 8'hf8;
    blue_mem[906] = 8'h1f;
    blue_mem[907] = 8'h80;
    blue_mem[908] = 8'hff;
    blue_mem[909] = 8'h7f;
    blue_mem[910] = 8'h00;
    blue_mem[911] = 8'h00;
    blue_mem[912] = 8'h00;
    blue_mem[913] = 8'h00;
    blue_mem[914] = 8'hfe;
    blue_mem[915] = 8'hff;
    blue_mem[916] = 8'hff;
    blue_mem[917] = 8'h1f;
    blue_mem[918] = 8'he0;
    blue_mem[919] = 8'hff;
    blue_mem[920] = 8'h03;
    blue_mem[921] = 8'hfe;
    blue_mem[922] = 8'h07;
    blue_mem[923] = 8'hf0;
    blue_mem[924] = 8'hff;
    blue_mem[925] = 8'h7f;
    blue_mem[926] = 8'h00;
    blue_mem[927] = 8'h00;
    blue_mem[928] = 8'h00;
    blue_mem[929] = 8'h00;
    blue_mem[930] = 8'hfc;
    blue_mem[931] = 8'hff;
    blue_mem[932] = 8'hff;
    blue_mem[933] = 8'h0f;
    blue_mem[934] = 8'he0;
    blue_mem[935] = 8'hff;
    blue_mem[936] = 8'h9f;
    blue_mem[937] = 8'hff;
    blue_mem[938] = 8'h07;
    blue_mem[939] = 8'hf0;
    blue_mem[940] = 8'hff;
    blue_mem[941] = 8'h7f;
    blue_mem[942] = 8'h00;
    blue_mem[943] = 8'h00;
    blue_mem[944] = 8'h00;
    blue_mem[945] = 8'h00;
    blue_mem[946] = 8'hfc;
    blue_mem[947] = 8'hff;
    blue_mem[948] = 8'hff;
    blue_mem[949] = 8'h0f;
    blue_mem[950] = 8'hf0;
    blue_mem[951] = 8'hff;
    blue_mem[952] = 8'hff;
    blue_mem[953] = 8'h7f;
    blue_mem[954] = 8'h00;
    blue_mem[955] = 8'hf8;
    blue_mem[956] = 8'hff;
    blue_mem[957] = 8'hff;
    blue_mem[958] = 8'h00;
    blue_mem[959] = 8'h00;
    blue_mem[960] = 8'h00;
    blue_mem[961] = 8'h00;
    blue_mem[962] = 8'hf0;
    blue_mem[963] = 8'hff;
    blue_mem[964] = 8'hff;
    blue_mem[965] = 8'h07;
    blue_mem[966] = 8'hf8;
    blue_mem[967] = 8'hff;
    blue_mem[968] = 8'hff;
    blue_mem[969] = 8'h7f;
    blue_mem[970] = 8'h00;
    blue_mem[971] = 8'hfc;
    blue_mem[972] = 8'hff;
    blue_mem[973] = 8'hff;
    blue_mem[974] = 8'h00;
    blue_mem[975] = 8'h00;
    blue_mem[976] = 8'h00;
    blue_mem[977] = 8'h00;
    blue_mem[978] = 8'hff;
    blue_mem[979] = 8'hff;
    blue_mem[980] = 8'hff;
    blue_mem[981] = 8'h0f;
    blue_mem[982] = 8'hf8;
    blue_mem[983] = 8'hff;
    blue_mem[984] = 8'hff;
    blue_mem[985] = 8'h77;
    blue_mem[986] = 8'h00;
    blue_mem[987] = 8'hff;
    blue_mem[988] = 8'hfd;
    blue_mem[989] = 8'h7f;
    blue_mem[990] = 8'h00;
    blue_mem[991] = 8'h00;
    blue_mem[992] = 8'h00;
    blue_mem[993] = 8'h00;
    blue_mem[994] = 8'hff;
    blue_mem[995] = 8'hff;
    blue_mem[996] = 8'hff;
    blue_mem[997] = 8'h0f;
    blue_mem[998] = 8'hf8;
    blue_mem[999] = 8'hff;
    blue_mem[1000] = 8'hff;
    blue_mem[1001] = 8'h7f;
    blue_mem[1002] = 8'h00;
    blue_mem[1003] = 8'hff;
    blue_mem[1004] = 8'hef;
    blue_mem[1005] = 8'h7f;
    blue_mem[1006] = 8'h00;
    blue_mem[1007] = 8'h00;
    blue_mem[1008] = 8'h00;
    blue_mem[1009] = 8'h00;
    blue_mem[1010] = 8'hff;
    blue_mem[1011] = 8'hff;
    blue_mem[1012] = 8'hff;
    blue_mem[1013] = 8'h0f;
    blue_mem[1014] = 8'hf8;
    blue_mem[1015] = 8'hff;
    blue_mem[1016] = 8'hff;
    blue_mem[1017] = 8'h1f;
    blue_mem[1018] = 8'he0;
    blue_mem[1019] = 8'hff;
    blue_mem[1020] = 8'hff;
    blue_mem[1021] = 8'h3f;
    blue_mem[1022] = 8'h00;
    blue_mem[1023] = 8'h00;
    blue_mem[1024] = 8'h00;
    blue_mem[1025] = 8'h00;
    blue_mem[1026] = 8'hfe;
    blue_mem[1027] = 8'hff;
    blue_mem[1028] = 8'hff;
    blue_mem[1029] = 8'h07;
    blue_mem[1030] = 8'h78;
    blue_mem[1031] = 8'hff;
    blue_mem[1032] = 8'hff;
    blue_mem[1033] = 8'h07;
    blue_mem[1034] = 8'hf0;
    blue_mem[1035] = 8'hff;
    blue_mem[1036] = 8'hff;
    blue_mem[1037] = 8'h7f;
    blue_mem[1038] = 8'h00;
    blue_mem[1039] = 8'h00;
    blue_mem[1040] = 8'h00;
    blue_mem[1041] = 8'h00;
    blue_mem[1042] = 8'hfe;
    blue_mem[1043] = 8'hff;
    blue_mem[1044] = 8'hff;
    blue_mem[1045] = 8'h07;
    blue_mem[1046] = 8'hf8;
    blue_mem[1047] = 8'hff;
    blue_mem[1048] = 8'hff;
    blue_mem[1049] = 8'h03;
    blue_mem[1050] = 8'hf6;
    blue_mem[1051] = 8'hff;
    blue_mem[1052] = 8'hff;
    blue_mem[1053] = 8'he7;
    blue_mem[1054] = 8'h00;
    blue_mem[1055] = 8'h00;
    blue_mem[1056] = 8'h00;
    blue_mem[1057] = 8'h00;
    blue_mem[1058] = 8'hfe;
    blue_mem[1059] = 8'hff;
    blue_mem[1060] = 8'hff;
    blue_mem[1061] = 8'h07;
    blue_mem[1062] = 8'hfc;
    blue_mem[1063] = 8'hff;
    blue_mem[1064] = 8'hff;
    blue_mem[1065] = 8'h41;
    blue_mem[1066] = 8'hff;
    blue_mem[1067] = 8'hff;
    blue_mem[1068] = 8'hff;
    blue_mem[1069] = 8'h7f;
    blue_mem[1070] = 8'h00;
    blue_mem[1071] = 8'h00;
    blue_mem[1072] = 8'h00;
    blue_mem[1073] = 8'h00;
    blue_mem[1074] = 8'hfe;
    blue_mem[1075] = 8'hbf;
    blue_mem[1076] = 8'hff;
    blue_mem[1077] = 8'h03;
    blue_mem[1078] = 8'hfe;
    blue_mem[1079] = 8'hff;
    blue_mem[1080] = 8'h7e;
    blue_mem[1081] = 8'he0;
    blue_mem[1082] = 8'hff;
    blue_mem[1083] = 8'hff;
    blue_mem[1084] = 8'hff;
    blue_mem[1085] = 8'h7f;
    blue_mem[1086] = 8'h00;
    blue_mem[1087] = 8'h00;
    blue_mem[1088] = 8'h00;
    blue_mem[1089] = 8'h00;
    blue_mem[1090] = 8'hfe;
    blue_mem[1091] = 8'hff;
    blue_mem[1092] = 8'hff;
    blue_mem[1093] = 8'h03;
    blue_mem[1094] = 8'hfe;
    blue_mem[1095] = 8'hff;
    blue_mem[1096] = 8'h3e;
    blue_mem[1097] = 8'he0;
    blue_mem[1098] = 8'hef;
    blue_mem[1099] = 8'hff;
    blue_mem[1100] = 8'hff;
    blue_mem[1101] = 8'hff;
    blue_mem[1102] = 8'h00;
    blue_mem[1103] = 8'h00;
    blue_mem[1104] = 8'h00;
    blue_mem[1105] = 8'h00;
    blue_mem[1106] = 8'hfc;
    blue_mem[1107] = 8'hff;
    blue_mem[1108] = 8'hf7;
    blue_mem[1109] = 8'h03;
    blue_mem[1110] = 8'hfe;
    blue_mem[1111] = 8'hff;
    blue_mem[1112] = 8'h1f;
    blue_mem[1113] = 8'h78;
    blue_mem[1114] = 8'hff;
    blue_mem[1115] = 8'hff;
    blue_mem[1116] = 8'hff;
    blue_mem[1117] = 8'h7f;
    blue_mem[1118] = 8'h00;
    blue_mem[1119] = 8'h00;
    blue_mem[1120] = 8'h00;
    blue_mem[1121] = 8'h00;
    blue_mem[1122] = 8'hfc;
    blue_mem[1123] = 8'hbf;
    blue_mem[1124] = 8'hff;
    blue_mem[1125] = 8'h03;
    blue_mem[1126] = 8'hff;
    blue_mem[1127] = 8'hff;
    blue_mem[1128] = 8'h07;
    blue_mem[1129] = 8'hfc;
    blue_mem[1130] = 8'hff;
    blue_mem[1131] = 8'hff;
    blue_mem[1132] = 8'hff;
    blue_mem[1133] = 8'h7f;
    blue_mem[1134] = 8'h00;
    blue_mem[1135] = 8'h00;
    blue_mem[1136] = 8'h00;
    blue_mem[1137] = 8'h00;
    blue_mem[1138] = 8'hfe;
    blue_mem[1139] = 8'hff;
    blue_mem[1140] = 8'hff;
    blue_mem[1141] = 8'h03;
    blue_mem[1142] = 8'hfe;
    blue_mem[1143] = 8'hff;
    blue_mem[1144] = 8'h87;
    blue_mem[1145] = 8'hff;
    blue_mem[1146] = 8'hff;
    blue_mem[1147] = 8'hff;
    blue_mem[1148] = 8'hff;
    blue_mem[1149] = 8'h7f;
    blue_mem[1150] = 8'h00;
    blue_mem[1151] = 8'h00;
    blue_mem[1152] = 8'h00;
    blue_mem[1153] = 8'h00;
    blue_mem[1154] = 8'hfe;
    blue_mem[1155] = 8'hff;
    blue_mem[1156] = 8'hff;
    blue_mem[1157] = 8'h01;
    blue_mem[1158] = 8'hfe;
    blue_mem[1159] = 8'hfb;
    blue_mem[1160] = 8'h80;
    blue_mem[1161] = 8'hff;
    blue_mem[1162] = 8'hff;
    blue_mem[1163] = 8'hff;
    blue_mem[1164] = 8'hff;
    blue_mem[1165] = 8'h7f;
    blue_mem[1166] = 8'h00;
    blue_mem[1167] = 8'h00;
    blue_mem[1168] = 8'h00;
    blue_mem[1169] = 8'h00;
    blue_mem[1170] = 8'hfc;
    blue_mem[1171] = 8'hff;
    blue_mem[1172] = 8'hff;
    blue_mem[1173] = 8'h03;
    blue_mem[1174] = 8'hfe;
    blue_mem[1175] = 8'h7f;
    blue_mem[1176] = 8'h00;
    blue_mem[1177] = 8'hfd;
    blue_mem[1178] = 8'hef;
    blue_mem[1179] = 8'hff;
    blue_mem[1180] = 8'hff;
    blue_mem[1181] = 8'h7e;
    blue_mem[1182] = 8'h00;
    blue_mem[1183] = 8'h00;
    blue_mem[1184] = 8'h00;
    blue_mem[1185] = 8'h00;
    blue_mem[1186] = 8'hfc;
    blue_mem[1187] = 8'hff;
    blue_mem[1188] = 8'hff;
    blue_mem[1189] = 8'h03;
    blue_mem[1190] = 8'hfe;
    blue_mem[1191] = 8'h7f;
    blue_mem[1192] = 8'h00;
    blue_mem[1193] = 8'hd8;
    blue_mem[1194] = 8'hef;
    blue_mem[1195] = 8'hc7;
    blue_mem[1196] = 8'hff;
    blue_mem[1197] = 8'h3f;
    blue_mem[1198] = 8'h00;
    blue_mem[1199] = 8'h00;
    blue_mem[1200] = 8'h00;
    blue_mem[1201] = 8'h00;
    blue_mem[1202] = 8'hf8;
    blue_mem[1203] = 8'h7f;
    blue_mem[1204] = 8'hcf;
    blue_mem[1205] = 8'h03;
    blue_mem[1206] = 8'hfe;
    blue_mem[1207] = 8'h7f;
    blue_mem[1208] = 8'h00;
    blue_mem[1209] = 8'h80;
    blue_mem[1210] = 8'hff;
    blue_mem[1211] = 8'hc3;
    blue_mem[1212] = 8'hff;
    blue_mem[1213] = 8'h37;
    blue_mem[1214] = 8'h00;
    blue_mem[1215] = 8'h00;
    blue_mem[1216] = 8'h00;
    blue_mem[1217] = 8'h00;
    blue_mem[1218] = 8'hf8;
    blue_mem[1219] = 8'hff;
    blue_mem[1220] = 8'hff;
    blue_mem[1221] = 8'h00;
    blue_mem[1222] = 8'hff;
    blue_mem[1223] = 8'h0f;
    blue_mem[1224] = 8'h00;
    blue_mem[1225] = 8'h00;
    blue_mem[1226] = 8'hf8;
    blue_mem[1227] = 8'hf1;
    blue_mem[1228] = 8'hff;
    blue_mem[1229] = 8'h3f;
    blue_mem[1230] = 8'h00;
    blue_mem[1231] = 8'h00;
    blue_mem[1232] = 8'h00;
    blue_mem[1233] = 8'h00;
    blue_mem[1234] = 8'hb8;
    blue_mem[1235] = 8'hff;
    blue_mem[1236] = 8'hff;
    blue_mem[1237] = 8'h80;
    blue_mem[1238] = 8'hff;
    blue_mem[1239] = 8'h07;
    blue_mem[1240] = 8'h00;
    blue_mem[1241] = 8'h00;
    blue_mem[1242] = 8'h10;
    blue_mem[1243] = 8'hf0;
    blue_mem[1244] = 8'hff;
    blue_mem[1245] = 8'h1f;
    blue_mem[1246] = 8'h00;
    blue_mem[1247] = 8'h00;
    blue_mem[1248] = 8'h00;
    blue_mem[1249] = 8'h00;
    blue_mem[1250] = 8'hf0;
    blue_mem[1251] = 8'hdf;
    blue_mem[1252] = 8'hff;
    blue_mem[1253] = 8'h80;
    blue_mem[1254] = 8'hff;
    blue_mem[1255] = 8'h07;
    blue_mem[1256] = 8'h00;
    blue_mem[1257] = 8'h00;
    blue_mem[1258] = 8'h00;
    blue_mem[1259] = 8'hf8;
    blue_mem[1260] = 8'hef;
    blue_mem[1261] = 8'h1f;
    blue_mem[1262] = 8'h00;
    blue_mem[1263] = 8'h00;
    blue_mem[1264] = 8'h00;
    blue_mem[1265] = 8'h00;
    blue_mem[1266] = 8'hf0;
    blue_mem[1267] = 8'hff;
    blue_mem[1268] = 8'hff;
    blue_mem[1269] = 8'h80;
    blue_mem[1270] = 8'hff;
    blue_mem[1271] = 8'h07;
    blue_mem[1272] = 8'h00;
    blue_mem[1273] = 8'h00;
    blue_mem[1274] = 8'h00;
    blue_mem[1275] = 8'hf8;
    blue_mem[1276] = 8'hff;
    blue_mem[1277] = 8'h1f;
    blue_mem[1278] = 8'h00;
    blue_mem[1279] = 8'h00;
    blue_mem[1280] = 8'h00;
    blue_mem[1281] = 8'h00;
    blue_mem[1282] = 8'hf0;
    blue_mem[1283] = 8'hff;
    blue_mem[1284] = 8'hff;
    blue_mem[1285] = 8'h00;
    blue_mem[1286] = 8'hff;
    blue_mem[1287] = 8'h03;
    blue_mem[1288] = 8'h18;
    blue_mem[1289] = 8'h00;
    blue_mem[1290] = 8'h00;
    blue_mem[1291] = 8'hf8;
    blue_mem[1292] = 8'hff;
    blue_mem[1293] = 8'h0f;
    blue_mem[1294] = 8'h00;
    blue_mem[1295] = 8'h00;
    blue_mem[1296] = 8'h00;
    blue_mem[1297] = 8'h00;
    blue_mem[1298] = 8'he0;
    blue_mem[1299] = 8'hff;
    blue_mem[1300] = 8'h27;
    blue_mem[1301] = 8'h00;
    blue_mem[1302] = 8'hf9;
    blue_mem[1303] = 8'h80;
    blue_mem[1304] = 8'hff;
    blue_mem[1305] = 8'h00;
    blue_mem[1306] = 8'h00;
    blue_mem[1307] = 8'hfc;
    blue_mem[1308] = 8'hff;
    blue_mem[1309] = 8'h0f;
    blue_mem[1310] = 8'h00;
    blue_mem[1311] = 8'h00;
    blue_mem[1312] = 8'h00;
    blue_mem[1313] = 8'h00;
    blue_mem[1314] = 8'he0;
    blue_mem[1315] = 8'hff;
    blue_mem[1316] = 8'h03;
    blue_mem[1317] = 8'h00;
    blue_mem[1318] = 8'hf0;
    blue_mem[1319] = 8'hf0;
    blue_mem[1320] = 8'hff;
    blue_mem[1321] = 8'h01;
    blue_mem[1322] = 8'h00;
    blue_mem[1323] = 8'hfe;
    blue_mem[1324] = 8'hdf;
    blue_mem[1325] = 8'h0f;
    blue_mem[1326] = 8'h00;
    blue_mem[1327] = 8'h00;
    blue_mem[1328] = 8'h00;
    blue_mem[1329] = 8'h00;
    blue_mem[1330] = 8'he0;
    blue_mem[1331] = 8'hff;
    blue_mem[1332] = 8'h03;
    blue_mem[1333] = 8'h00;
    blue_mem[1334] = 8'hf0;
    blue_mem[1335] = 8'hf0;
    blue_mem[1336] = 8'hff;
    blue_mem[1337] = 8'h0f;
    blue_mem[1338] = 8'hc0;
    blue_mem[1339] = 8'hff;
    blue_mem[1340] = 8'hff;
    blue_mem[1341] = 8'h07;
    blue_mem[1342] = 8'h00;
    blue_mem[1343] = 8'h00;
    blue_mem[1344] = 8'h00;
    blue_mem[1345] = 8'h00;
    blue_mem[1346] = 8'h80;
    blue_mem[1347] = 8'hff;
    blue_mem[1348] = 8'h03;
    blue_mem[1349] = 8'h86;
    blue_mem[1350] = 8'hf0;
    blue_mem[1351] = 8'hf9;
    blue_mem[1352] = 8'hff;
    blue_mem[1353] = 8'hff;
    blue_mem[1354] = 8'hf8;
    blue_mem[1355] = 8'hff;
    blue_mem[1356] = 8'hff;
    blue_mem[1357] = 8'h07;
    blue_mem[1358] = 8'h00;
    blue_mem[1359] = 8'h00;
    blue_mem[1360] = 8'h00;
    blue_mem[1361] = 8'h00;
    blue_mem[1362] = 8'h80;
    blue_mem[1363] = 8'hff;
    blue_mem[1364] = 8'hf7;
    blue_mem[1365] = 8'hc7;
    blue_mem[1366] = 8'hfd;
    blue_mem[1367] = 8'hff;
    blue_mem[1368] = 8'hff;
    blue_mem[1369] = 8'hff;
    blue_mem[1370] = 8'hff;
    blue_mem[1371] = 8'hff;
    blue_mem[1372] = 8'hff;
    blue_mem[1373] = 8'h07;
    blue_mem[1374] = 8'h00;
    blue_mem[1375] = 8'h00;
    blue_mem[1376] = 8'h00;
    blue_mem[1377] = 8'h00;
    blue_mem[1378] = 8'hc0;
    blue_mem[1379] = 8'hff;
    blue_mem[1380] = 8'hff;
    blue_mem[1381] = 8'hff;
    blue_mem[1382] = 8'hfd;
    blue_mem[1383] = 8'hf7;
    blue_mem[1384] = 8'hff;
    blue_mem[1385] = 8'hff;
    blue_mem[1386] = 8'hff;
    blue_mem[1387] = 8'hff;
    blue_mem[1388] = 8'hff;
    blue_mem[1389] = 8'h07;
    blue_mem[1390] = 8'h00;
    blue_mem[1391] = 8'h00;
    blue_mem[1392] = 8'h00;
    blue_mem[1393] = 8'h00;
    blue_mem[1394] = 8'h00;
    blue_mem[1395] = 8'hff;
    blue_mem[1396] = 8'hff;
    blue_mem[1397] = 8'hfd;
    blue_mem[1398] = 8'hff;
    blue_mem[1399] = 8'hf7;
    blue_mem[1400] = 8'hff;
    blue_mem[1401] = 8'hff;
    blue_mem[1402] = 8'hff;
    blue_mem[1403] = 8'hff;
    blue_mem[1404] = 8'hff;
    blue_mem[1405] = 8'h03;
    blue_mem[1406] = 8'h00;
    blue_mem[1407] = 8'h00;
    blue_mem[1408] = 8'h00;
    blue_mem[1409] = 8'h00;
    blue_mem[1410] = 8'h00;
    blue_mem[1411] = 8'hff;
    blue_mem[1412] = 8'hff;
    blue_mem[1413] = 8'hff;
    blue_mem[1414] = 8'hff;
    blue_mem[1415] = 8'hff;
    blue_mem[1416] = 8'hff;
    blue_mem[1417] = 8'hff;
    blue_mem[1418] = 8'hf7;
    blue_mem[1419] = 8'hff;
    blue_mem[1420] = 8'hff;
    blue_mem[1421] = 8'h00;
    blue_mem[1422] = 8'h00;
    blue_mem[1423] = 8'h00;
    blue_mem[1424] = 8'h00;
    blue_mem[1425] = 8'h00;
    blue_mem[1426] = 8'h00;
    blue_mem[1427] = 8'hff;
    blue_mem[1428] = 8'hfe;
    blue_mem[1429] = 8'hf7;
    blue_mem[1430] = 8'hff;
    blue_mem[1431] = 8'hff;
    blue_mem[1432] = 8'hff;
    blue_mem[1433] = 8'hff;
    blue_mem[1434] = 8'hff;
    blue_mem[1435] = 8'hff;
    blue_mem[1436] = 8'hff;
    blue_mem[1437] = 8'h00;
    blue_mem[1438] = 8'h00;
    blue_mem[1439] = 8'h00;
    blue_mem[1440] = 8'h00;
    blue_mem[1441] = 8'h00;
    blue_mem[1442] = 8'h00;
    blue_mem[1443] = 8'hfc;
    blue_mem[1444] = 8'hef;
    blue_mem[1445] = 8'hff;
    blue_mem[1446] = 8'hff;
    blue_mem[1447] = 8'hff;
    blue_mem[1448] = 8'hff;
    blue_mem[1449] = 8'hff;
    blue_mem[1450] = 8'hff;
    blue_mem[1451] = 8'hff;
    blue_mem[1452] = 8'hff;
    blue_mem[1453] = 8'h00;
    blue_mem[1454] = 8'h00;
    blue_mem[1455] = 8'h00;
    blue_mem[1456] = 8'h00;
    blue_mem[1457] = 8'h00;
    blue_mem[1458] = 8'h00;
    blue_mem[1459] = 8'hfc;
    blue_mem[1460] = 8'hff;
    blue_mem[1461] = 8'hff;
    blue_mem[1462] = 8'hff;
    blue_mem[1463] = 8'hff;
    blue_mem[1464] = 8'h9f;
    blue_mem[1465] = 8'hff;
    blue_mem[1466] = 8'hff;
    blue_mem[1467] = 8'hff;
    blue_mem[1468] = 8'h3f;
    blue_mem[1469] = 8'h00;
    blue_mem[1470] = 8'h00;
    blue_mem[1471] = 8'h00;
    blue_mem[1472] = 8'h00;
    blue_mem[1473] = 8'h00;
    blue_mem[1474] = 8'h00;
    blue_mem[1475] = 8'hf8;
    blue_mem[1476] = 8'hff;
    blue_mem[1477] = 8'hff;
    blue_mem[1478] = 8'hff;
    blue_mem[1479] = 8'hff;
    blue_mem[1480] = 8'hff;
    blue_mem[1481] = 8'hff;
    blue_mem[1482] = 8'hff;
    blue_mem[1483] = 8'hff;
    blue_mem[1484] = 8'h3f;
    blue_mem[1485] = 8'h00;
    blue_mem[1486] = 8'h00;
    blue_mem[1487] = 8'h00;
    blue_mem[1488] = 8'h00;
    blue_mem[1489] = 8'h00;
    blue_mem[1490] = 8'h00;
    blue_mem[1491] = 8'h70;
    blue_mem[1492] = 8'h7f;
    blue_mem[1493] = 8'hff;
    blue_mem[1494] = 8'hff;
    blue_mem[1495] = 8'hff;
    blue_mem[1496] = 8'hf7;
    blue_mem[1497] = 8'hff;
    blue_mem[1498] = 8'hff;
    blue_mem[1499] = 8'hf7;
    blue_mem[1500] = 8'h1f;
    blue_mem[1501] = 8'h00;
    blue_mem[1502] = 8'h00;
    blue_mem[1503] = 8'h00;
    blue_mem[1504] = 8'h00;
    blue_mem[1505] = 8'h00;
    blue_mem[1506] = 8'h00;
    blue_mem[1507] = 8'he0;
    blue_mem[1508] = 8'hff;
    blue_mem[1509] = 8'hff;
    blue_mem[1510] = 8'hff;
    blue_mem[1511] = 8'hff;
    blue_mem[1512] = 8'hf7;
    blue_mem[1513] = 8'hef;
    blue_mem[1514] = 8'hff;
    blue_mem[1515] = 8'hff;
    blue_mem[1516] = 8'h0f;
    blue_mem[1517] = 8'h00;
    blue_mem[1518] = 8'h00;
    blue_mem[1519] = 8'h00;
    blue_mem[1520] = 8'h00;
    blue_mem[1521] = 8'h00;
    blue_mem[1522] = 8'h00;
    blue_mem[1523] = 8'he0;
    blue_mem[1524] = 8'hfd;
    blue_mem[1525] = 8'hff;
    blue_mem[1526] = 8'hff;
    blue_mem[1527] = 8'hff;
    blue_mem[1528] = 8'hff;
    blue_mem[1529] = 8'hff;
    blue_mem[1530] = 8'hff;
    blue_mem[1531] = 8'hff;
    blue_mem[1532] = 8'h03;
    blue_mem[1533] = 8'h00;
    blue_mem[1534] = 8'h00;
    blue_mem[1535] = 8'h00;
    blue_mem[1536] = 8'h00;
    blue_mem[1537] = 8'h00;
    blue_mem[1538] = 8'h00;
    blue_mem[1539] = 8'hc0;
    blue_mem[1540] = 8'hff;
    blue_mem[1541] = 8'hff;
    blue_mem[1542] = 8'hff;
    blue_mem[1543] = 8'hef;
    blue_mem[1544] = 8'hff;
    blue_mem[1545] = 8'hff;
    blue_mem[1546] = 8'h7b;
    blue_mem[1547] = 8'hff;
    blue_mem[1548] = 8'h01;
    blue_mem[1549] = 8'h00;
    blue_mem[1550] = 8'h00;
    blue_mem[1551] = 8'h00;
    blue_mem[1552] = 8'h00;
    blue_mem[1553] = 8'h00;
    blue_mem[1554] = 8'h00;
    blue_mem[1555] = 8'h00;
    blue_mem[1556] = 8'hff;
    blue_mem[1557] = 8'hff;
    blue_mem[1558] = 8'hff;
    blue_mem[1559] = 8'hff;
    blue_mem[1560] = 8'hff;
    blue_mem[1561] = 8'hff;
    blue_mem[1562] = 8'hff;
    blue_mem[1563] = 8'hff;
    blue_mem[1564] = 8'h00;
    blue_mem[1565] = 8'h00;
    blue_mem[1566] = 8'h00;
    blue_mem[1567] = 8'h00;
    blue_mem[1568] = 8'h00;
    blue_mem[1569] = 8'h00;
    blue_mem[1570] = 8'h00;
    blue_mem[1571] = 8'h00;
    blue_mem[1572] = 8'hef;
    blue_mem[1573] = 8'hff;
    blue_mem[1574] = 8'hff;
    blue_mem[1575] = 8'hff;
    blue_mem[1576] = 8'hff;
    blue_mem[1577] = 8'hff;
    blue_mem[1578] = 8'hff;
    blue_mem[1579] = 8'hff;
    blue_mem[1580] = 8'h00;
    blue_mem[1581] = 8'h00;
    blue_mem[1582] = 8'h00;
    blue_mem[1583] = 8'h00;
    blue_mem[1584] = 8'h00;
    blue_mem[1585] = 8'h00;
    blue_mem[1586] = 8'h00;
    blue_mem[1587] = 8'h00;
    blue_mem[1588] = 8'hfe;
    blue_mem[1589] = 8'hff;
    blue_mem[1590] = 8'hff;
    blue_mem[1591] = 8'hff;
    blue_mem[1592] = 8'hff;
    blue_mem[1593] = 8'hff;
    blue_mem[1594] = 8'hff;
    blue_mem[1595] = 8'h7f;
    blue_mem[1596] = 8'h00;
    blue_mem[1597] = 8'h00;
    blue_mem[1598] = 8'h00;
    blue_mem[1599] = 8'h00;
    blue_mem[1600] = 8'h00;
    blue_mem[1601] = 8'h00;
    blue_mem[1602] = 8'h00;
    blue_mem[1603] = 8'h00;
    blue_mem[1604] = 8'hf0;
    blue_mem[1605] = 8'hff;
    blue_mem[1606] = 8'hff;
    blue_mem[1607] = 8'hff;
    blue_mem[1608] = 8'hff;
    blue_mem[1609] = 8'hff;
    blue_mem[1610] = 8'hff;
    blue_mem[1611] = 8'h1f;
    blue_mem[1612] = 8'h00;
    blue_mem[1613] = 8'h00;
    blue_mem[1614] = 8'h00;
    blue_mem[1615] = 8'h00;
    blue_mem[1616] = 8'h00;
    blue_mem[1617] = 8'h00;
    blue_mem[1618] = 8'h00;
    blue_mem[1619] = 8'h00;
    blue_mem[1620] = 8'hf0;
    blue_mem[1621] = 8'hff;
    blue_mem[1622] = 8'hff;
    blue_mem[1623] = 8'hff;
    blue_mem[1624] = 8'hf7;
    blue_mem[1625] = 8'hff;
    blue_mem[1626] = 8'hff;
    blue_mem[1627] = 8'h1f;
    blue_mem[1628] = 8'h00;
    blue_mem[1629] = 8'h00;
    blue_mem[1630] = 8'h00;
    blue_mem[1631] = 8'h00;
    blue_mem[1632] = 8'h00;
    blue_mem[1633] = 8'h00;
    blue_mem[1634] = 8'h00;
    blue_mem[1635] = 8'h00;
    blue_mem[1636] = 8'he0;
    blue_mem[1637] = 8'hff;
    blue_mem[1638] = 8'hf6;
    blue_mem[1639] = 8'hef;
    blue_mem[1640] = 8'hff;
    blue_mem[1641] = 8'hfd;
    blue_mem[1642] = 8'hff;
    blue_mem[1643] = 8'h07;
    blue_mem[1644] = 8'h00;
    blue_mem[1645] = 8'h00;
    blue_mem[1646] = 8'h00;
    blue_mem[1647] = 8'h00;
    blue_mem[1648] = 8'h00;
    blue_mem[1649] = 8'h00;
    blue_mem[1650] = 8'h00;
    blue_mem[1651] = 8'h00;
    blue_mem[1652] = 8'h00;
    blue_mem[1653] = 8'h7e;
    blue_mem[1654] = 8'hff;
    blue_mem[1655] = 8'hff;
    blue_mem[1656] = 8'hff;
    blue_mem[1657] = 8'hff;
    blue_mem[1658] = 8'hff;
    blue_mem[1659] = 8'h03;
    blue_mem[1660] = 8'h00;
    blue_mem[1661] = 8'h00;
    blue_mem[1662] = 8'h00;
    blue_mem[1663] = 8'h00;
    blue_mem[1664] = 8'h00;
    blue_mem[1665] = 8'h00;
    blue_mem[1666] = 8'h00;
    blue_mem[1667] = 8'h00;
    blue_mem[1668] = 8'h00;
    blue_mem[1669] = 8'hfe;
    blue_mem[1670] = 8'hff;
    blue_mem[1671] = 8'hff;
    blue_mem[1672] = 8'hcf;
    blue_mem[1673] = 8'hff;
    blue_mem[1674] = 8'hff;
    blue_mem[1675] = 8'h00;
    blue_mem[1676] = 8'h00;
    blue_mem[1677] = 8'h00;
    blue_mem[1678] = 8'h00;
    blue_mem[1679] = 8'h00;
    blue_mem[1680] = 8'h00;
    blue_mem[1681] = 8'h00;
    blue_mem[1682] = 8'h00;
    blue_mem[1683] = 8'h00;
    blue_mem[1684] = 8'h00;
    blue_mem[1685] = 8'hf8;
    blue_mem[1686] = 8'hff;
    blue_mem[1687] = 8'hdf;
    blue_mem[1688] = 8'hff;
    blue_mem[1689] = 8'hfc;
    blue_mem[1690] = 8'h3f;
    blue_mem[1691] = 8'h00;
    blue_mem[1692] = 8'h00;
    blue_mem[1693] = 8'h00;
    blue_mem[1694] = 8'h00;
    blue_mem[1695] = 8'h00;
    blue_mem[1696] = 8'h00;
    blue_mem[1697] = 8'h00;
    blue_mem[1698] = 8'h00;
    blue_mem[1699] = 8'h00;
    blue_mem[1700] = 8'h00;
    blue_mem[1701] = 8'hf0;
    blue_mem[1702] = 8'hff;
    blue_mem[1703] = 8'hff;
    blue_mem[1704] = 8'hfb;
    blue_mem[1705] = 8'hff;
    blue_mem[1706] = 8'h1f;
    blue_mem[1707] = 8'h00;
    blue_mem[1708] = 8'h00;
    blue_mem[1709] = 8'h00;
    blue_mem[1710] = 8'h00;
    blue_mem[1711] = 8'h00;
    blue_mem[1712] = 8'h00;
    blue_mem[1713] = 8'h00;
    blue_mem[1714] = 8'h00;
    blue_mem[1715] = 8'h00;
    blue_mem[1716] = 8'h00;
    blue_mem[1717] = 8'h00;
    blue_mem[1718] = 8'hff;
    blue_mem[1719] = 8'hff;
    blue_mem[1720] = 8'hff;
    blue_mem[1721] = 8'hff;
    blue_mem[1722] = 8'h01;
    blue_mem[1723] = 8'h00;
    blue_mem[1724] = 8'h00;
    blue_mem[1725] = 8'h00;
    blue_mem[1726] = 8'h00;
    blue_mem[1727] = 8'h00;
    blue_mem[1728] = 8'h00;
    blue_mem[1729] = 8'h00;
    blue_mem[1730] = 8'h00;
    blue_mem[1731] = 8'h00;
    blue_mem[1732] = 8'h00;
    blue_mem[1733] = 8'h00;
    blue_mem[1734] = 8'hfe;
    blue_mem[1735] = 8'hff;
    blue_mem[1736] = 8'hff;
    blue_mem[1737] = 8'h3f;
    blue_mem[1738] = 8'h00;
    blue_mem[1739] = 8'h00;
    blue_mem[1740] = 8'h00;
    blue_mem[1741] = 8'h00;
    blue_mem[1742] = 8'h00;
    blue_mem[1743] = 8'h00;
    blue_mem[1744] = 8'h00;
    blue_mem[1745] = 8'h00;
    blue_mem[1746] = 8'h00;
    blue_mem[1747] = 8'h00;
    blue_mem[1748] = 8'h00;
    blue_mem[1749] = 8'h00;
    blue_mem[1750] = 8'h18;
    blue_mem[1751] = 8'hfe;
    blue_mem[1752] = 8'hff;
    blue_mem[1753] = 8'h1f;
    blue_mem[1754] = 8'h00;
    blue_mem[1755] = 8'h00;
    blue_mem[1756] = 8'h00;
    blue_mem[1757] = 8'h00;
    blue_mem[1758] = 8'h00;
    blue_mem[1759] = 8'h00;
    blue_mem[1760] = 8'h00;
    blue_mem[1761] = 8'h00;
    blue_mem[1762] = 8'h00;
    blue_mem[1763] = 8'h00;
    blue_mem[1764] = 8'h00;
    blue_mem[1765] = 8'h00;
    blue_mem[1766] = 8'h00;
    blue_mem[1767] = 8'hee;
    blue_mem[1768] = 8'hff;
    blue_mem[1769] = 8'h00;
    blue_mem[1770] = 8'h00;
    blue_mem[1771] = 8'h00;
    blue_mem[1772] = 8'h00;
    blue_mem[1773] = 8'h00;
    blue_mem[1774] = 8'h00;
    blue_mem[1775] = 8'h00;
    blue_mem[1776] = 8'h00;
    blue_mem[1777] = 8'h00;
    blue_mem[1778] = 8'h00;
    blue_mem[1779] = 8'h00;
    blue_mem[1780] = 8'h00;
    blue_mem[1781] = 8'h00;
    blue_mem[1782] = 8'h00;
    blue_mem[1783] = 8'h00;
    blue_mem[1784] = 8'h0c;
    blue_mem[1785] = 8'h00;
    blue_mem[1786] = 8'h00;
    blue_mem[1787] = 8'h00;
    blue_mem[1788] = 8'h00;
    blue_mem[1789] = 8'h00;
    blue_mem[1790] = 8'h00;
    blue_mem[1791] = 8'h00;
    blue_mem[1792] = 8'h00;
    blue_mem[1793] = 8'h00;
    blue_mem[1794] = 8'h00;
    blue_mem[1795] = 8'h00;
    blue_mem[1796] = 8'h00;
    blue_mem[1797] = 8'h00;
    blue_mem[1798] = 8'h00;
    blue_mem[1799] = 8'h00;
    blue_mem[1800] = 8'h00;
    blue_mem[1801] = 8'h00;
    blue_mem[1802] = 8'h00;
    blue_mem[1803] = 8'h00;
    blue_mem[1804] = 8'h00;
    blue_mem[1805] = 8'h00;
    blue_mem[1806] = 8'h00;
    blue_mem[1807] = 8'h00;
    blue_mem[1808] = 8'h00;
    blue_mem[1809] = 8'h00;
    blue_mem[1810] = 8'h00;
    blue_mem[1811] = 8'h00;
    blue_mem[1812] = 8'h00;
    blue_mem[1813] = 8'h00;
    blue_mem[1814] = 8'h00;
    blue_mem[1815] = 8'h00;
    blue_mem[1816] = 8'h00;
    blue_mem[1817] = 8'h00;
    blue_mem[1818] = 8'h00;
    blue_mem[1819] = 8'h00;
    blue_mem[1820] = 8'h00;
    blue_mem[1821] = 8'h00;
    blue_mem[1822] = 8'h00;
    blue_mem[1823] = 8'h00;
    blue_mem[1824] = 8'h00;
    blue_mem[1825] = 8'h00;
    blue_mem[1826] = 8'h00;
    blue_mem[1827] = 8'h00;
    blue_mem[1828] = 8'h00;
    blue_mem[1829] = 8'h00;
    blue_mem[1830] = 8'h00;
    blue_mem[1831] = 8'h00;
    blue_mem[1832] = 8'h00;
    blue_mem[1833] = 8'h00;
    blue_mem[1834] = 8'h00;
    blue_mem[1835] = 8'h00;
    blue_mem[1836] = 8'h00;
    blue_mem[1837] = 8'h00;
    blue_mem[1838] = 8'h00;
    blue_mem[1839] = 8'h00;
    blue_mem[1840] = 8'h00;
    blue_mem[1841] = 8'h00;
    blue_mem[1842] = 8'h00;
    blue_mem[1843] = 8'h00;
    blue_mem[1844] = 8'h00;
    blue_mem[1845] = 8'h00;
    blue_mem[1846] = 8'h00;
    blue_mem[1847] = 8'h00;
    blue_mem[1848] = 8'h00;
    blue_mem[1849] = 8'h00;
    blue_mem[1850] = 8'h00;
    blue_mem[1851] = 8'h00;
    blue_mem[1852] = 8'h00;
    blue_mem[1853] = 8'h00;
    blue_mem[1854] = 8'h00;
    blue_mem[1855] = 8'h00;
    blue_mem[1856] = 8'h00;
    blue_mem[1857] = 8'h00;
    blue_mem[1858] = 8'h00;
    blue_mem[1859] = 8'h00;
    blue_mem[1860] = 8'h00;
    blue_mem[1861] = 8'h00;
    blue_mem[1862] = 8'h00;
    blue_mem[1863] = 8'h00;
    blue_mem[1864] = 8'h00;
    blue_mem[1865] = 8'h00;
    blue_mem[1866] = 8'h00;
    blue_mem[1867] = 8'h00;
    blue_mem[1868] = 8'h00;
    blue_mem[1869] = 8'h00;
    blue_mem[1870] = 8'h00;
    blue_mem[1871] = 8'h00;
    blue_mem[1872] = 8'h00;
    blue_mem[1873] = 8'h00;
    blue_mem[1874] = 8'h00;
    blue_mem[1875] = 8'h00;
    blue_mem[1876] = 8'h00;
    blue_mem[1877] = 8'h00;
    blue_mem[1878] = 8'h00;
    blue_mem[1879] = 8'h00;
    blue_mem[1880] = 8'h00;
    blue_mem[1881] = 8'h00;
    blue_mem[1882] = 8'h00;
    blue_mem[1883] = 8'h00;
    blue_mem[1884] = 8'h00;
    blue_mem[1885] = 8'h00;
    blue_mem[1886] = 8'h00;
    blue_mem[1887] = 8'h00;
    blue_mem[1888] = 8'h00;
    blue_mem[1889] = 8'h00;
    blue_mem[1890] = 8'h00;
    blue_mem[1891] = 8'h00;
    blue_mem[1892] = 8'h00;
    blue_mem[1893] = 8'h00;
    blue_mem[1894] = 8'h00;
    blue_mem[1895] = 8'h00;
    blue_mem[1896] = 8'h00;
    blue_mem[1897] = 8'h00;
    blue_mem[1898] = 8'h00;
    blue_mem[1899] = 8'h00;
    blue_mem[1900] = 8'h00;
    blue_mem[1901] = 8'h00;
    blue_mem[1902] = 8'h00;
    blue_mem[1903] = 8'h00;
    blue_mem[1904] = 8'h00;
    blue_mem[1905] = 8'h00;
    blue_mem[1906] = 8'h00;
    blue_mem[1907] = 8'h00;
    blue_mem[1908] = 8'h00;
    blue_mem[1909] = 8'h00;
    blue_mem[1910] = 8'h00;
    blue_mem[1911] = 8'h00;
    blue_mem[1912] = 8'h00;
    blue_mem[1913] = 8'h00;
    blue_mem[1914] = 8'h00;
    blue_mem[1915] = 8'h00;
    blue_mem[1916] = 8'h00;
    blue_mem[1917] = 8'h00;
    blue_mem[1918] = 8'h00;
    blue_mem[1919] = 8'h00;
    blue_mem[1920] = 8'h00;
    blue_mem[1921] = 8'h00;
    blue_mem[1922] = 8'h00;
    blue_mem[1923] = 8'h00;
    blue_mem[1924] = 8'h00;
    blue_mem[1925] = 8'h00;
    blue_mem[1926] = 8'h00;
    blue_mem[1927] = 8'h00;
    blue_mem[1928] = 8'h00;
    blue_mem[1929] = 8'h00;
    blue_mem[1930] = 8'h00;
    blue_mem[1931] = 8'h00;
    blue_mem[1932] = 8'h00;
    blue_mem[1933] = 8'h00;
    blue_mem[1934] = 8'h00;
    blue_mem[1935] = 8'h00;
    blue_mem[1936] = 8'h00;
    blue_mem[1937] = 8'h00;
    blue_mem[1938] = 8'h00;
    blue_mem[1939] = 8'h00;
    blue_mem[1940] = 8'h00;
    blue_mem[1941] = 8'h00;
    blue_mem[1942] = 8'h00;
    blue_mem[1943] = 8'h00;
    blue_mem[1944] = 8'h00;
    blue_mem[1945] = 8'h00;
    blue_mem[1946] = 8'h00;
    blue_mem[1947] = 8'h00;
    blue_mem[1948] = 8'h00;
    blue_mem[1949] = 8'h00;
    blue_mem[1950] = 8'h00;
    blue_mem[1951] = 8'h00;
    blue_mem[1952] = 8'h00;
    blue_mem[1953] = 8'h00;
    blue_mem[1954] = 8'h00;
    blue_mem[1955] = 8'h00;
    blue_mem[1956] = 8'h00;
    blue_mem[1957] = 8'h00;
    blue_mem[1958] = 8'h00;
    blue_mem[1959] = 8'h00;
    blue_mem[1960] = 8'h00;
    blue_mem[1961] = 8'h00;
    blue_mem[1962] = 8'h00;
    blue_mem[1963] = 8'h00;
    blue_mem[1964] = 8'h00;
    blue_mem[1965] = 8'h00;
    blue_mem[1966] = 8'h00;
    blue_mem[1967] = 8'h00;
    blue_mem[1968] = 8'h00;
    blue_mem[1969] = 8'h00;
    blue_mem[1970] = 8'h00;
    blue_mem[1971] = 8'h00;
    blue_mem[1972] = 8'h00;
    blue_mem[1973] = 8'h00;
    blue_mem[1974] = 8'h00;
    blue_mem[1975] = 8'h00;
    blue_mem[1976] = 8'h00;
    blue_mem[1977] = 8'h00;
    blue_mem[1978] = 8'h00;
    blue_mem[1979] = 8'h00;
    blue_mem[1980] = 8'h00;
    blue_mem[1981] = 8'h00;
    blue_mem[1982] = 8'h00;
    blue_mem[1983] = 8'h00;
    blue_mem[1984] = 8'h00;
    blue_mem[1985] = 8'h00;
    blue_mem[1986] = 8'h00;
    blue_mem[1987] = 8'h00;
    blue_mem[1988] = 8'h00;
    blue_mem[1989] = 8'h00;
    blue_mem[1990] = 8'h00;
    blue_mem[1991] = 8'h00;
    blue_mem[1992] = 8'h00;
    blue_mem[1993] = 8'h00;
    blue_mem[1994] = 8'h00;
    blue_mem[1995] = 8'h00;
    blue_mem[1996] = 8'h00;
    blue_mem[1997] = 8'h00;
    blue_mem[1998] = 8'h00;
    blue_mem[1999] = 8'h00;
    blue_mem[2000] = 8'h00;
    blue_mem[2001] = 8'h00;
    blue_mem[2002] = 8'h00;
    blue_mem[2003] = 8'h00;
    blue_mem[2004] = 8'h00;
    blue_mem[2005] = 8'h00;
    blue_mem[2006] = 8'h00;
    blue_mem[2007] = 8'h00;
    blue_mem[2008] = 8'h00;
    blue_mem[2009] = 8'h00;
    blue_mem[2010] = 8'h00;
    blue_mem[2011] = 8'h00;
    blue_mem[2012] = 8'h00;
    blue_mem[2013] = 8'h00;
    blue_mem[2014] = 8'h00;
    blue_mem[2015] = 8'h00;
    blue_mem[2016] = 8'h00;
    blue_mem[2017] = 8'h00;
    blue_mem[2018] = 8'h00;
    blue_mem[2019] = 8'h00;
    blue_mem[2020] = 8'h00;
    blue_mem[2021] = 8'h00;
    blue_mem[2022] = 8'h00;
    blue_mem[2023] = 8'h00;
    blue_mem[2024] = 8'h00;
    blue_mem[2025] = 8'h00;
    blue_mem[2026] = 8'h00;
    blue_mem[2027] = 8'h00;
    blue_mem[2028] = 8'h00;
    blue_mem[2029] = 8'h00;
    blue_mem[2030] = 8'h00;
    blue_mem[2031] = 8'h00;
    blue_mem[2032] = 8'h00;
    blue_mem[2033] = 8'h00;
    blue_mem[2034] = 8'h00;
    blue_mem[2035] = 8'h00;
    blue_mem[2036] = 8'h00;
    blue_mem[2037] = 8'h00;
    blue_mem[2038] = 8'h00;
    blue_mem[2039] = 8'h00;
    blue_mem[2040] = 8'h00;
    blue_mem[2041] = 8'h00;
    blue_mem[2042] = 8'h00;
    blue_mem[2043] = 8'h00;
    blue_mem[2044] = 8'h00;
    blue_mem[2045] = 8'h00;
    blue_mem[2046] = 8'h00;
    blue_mem[2047] = 8'h00;
  end

  wire [10:0] addr = {y[6:0], x[6:3]};
  assign red_pixel = red_mem[addr][x&7];
  assign green_pixel = green_mem[addr][x&7];
  assign blue_pixel = blue_mem[addr][x&7];

endmodule

/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none
`define COLOR_WHITE 3'd7

module tt_um_vga_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // VGA signals
  wire hsync;
  wire vsync;
  reg [1:0] R;
  reg [1:0] G;
  reg [1:0] B;
  wire video_active;
  wire [9:0] pix_x;
  wire [9:0] pix_y;

  // Configuration
  wire cfg_tile = ui_in[0];
  wire cfg_solid_color = ui_in[1];

  // TinyVGA PMOD
  assign uo_out  = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};

  // Unused outputs assigned to 0.
  assign uio_out = 0;
  assign uio_oe  = 0;

  // Suppress unused signals warning
  wire _unused_ok = &{ena, ui_in[7:1], uio_in};

  vga_sync_generator vga_sync_gen (
      .clk(clk),
      .reset(~rst_n),
      .hsync(hsync),
      .vsync(vsync),
      .display_on(video_active),
      .hpos(pix_x),
      .vpos(pix_y)
  );


  wire pixel_value;
  wire [5:0] pallete_color;
  wire [5:0] color;

  wire [9:0] x = pix_x - logo_left;
  wire [9:0] y = pix_y - logo_top;
  wire logo_pixels = cfg_tile || (x[9:7] == 0 && y[9:7] == 0);

  bitmap_rom rom1 (
      .x(x[6:0]),
      .y(y[6:0]),
      .pixel(pixel_value)
  );

  palette palette_inst (
      .color_index(color_index),
      .rrggbb(pallete_color)
  );

  wire [5:0] gradient_color = {1'b1, y[6:2] - x[6:2] + logo_left[6:2]};
  assign color = cfg_solid_color ? pallete_color : gradient_color;

  // RGB output logic
  always @(posedge clk) begin
    if (~rst_n) begin
      R <= 0;
      G <= 0;
      B <= 0;
    end else begin
      R <= 0;
      G <= 0;
      B <= 0;
      if (video_active && logo_pixels) begin
        R <= pixel_value ? color[5:4] : 0;
        G <= pixel_value ? color[3:2] : 0;
        B <= pixel_value ? color[1:0] : 0;
      end
    end
  end

endmodule

module bitmap_rom (
    input wire [6:0] x,
    input wire [6:1] y,
    output wire pixel
);

  reg [5:0] mem[4095:0];
  initial begin

mem[0] = 6'b111111;
mem[1] = 6'b111111;
mem[2] = 6'b111111;
mem[3] = 6'b111111;
mem[4] = 6'b111111;
mem[5] = 6'b111111;
mem[6] = 6'b111111;
mem[7] = 6'b111111;
mem[8] = 6'b111111;
mem[9] = 6'b111111;
mem[10] = 6'b111111;
mem[11] = 6'b111111;
mem[12] = 6'b111111;
mem[13] = 6'b111111;
mem[14] = 6'b111111;
mem[15] = 6'b111111;
mem[16] = 6'b111111;
mem[17] = 6'b111111;
mem[18] = 6'b111111;
mem[19] = 6'b111111;
mem[20] = 6'b111111;
mem[21] = 6'b111111;
mem[22] = 6'b111111;
mem[23] = 6'b111111;
mem[24] = 6'b111111;
mem[25] = 6'b111111;
mem[26] = 6'b111111;
mem[27] = 6'b111111;
mem[28] = 6'b111111;
mem[29] = 6'b111111;
mem[30] = 6'b111111;
mem[31] = 6'b111111;
mem[32] = 6'b111111;
mem[33] = 6'b111111;
mem[34] = 6'b111111;
mem[35] = 6'b111111;
mem[36] = 6'b111111;
mem[37] = 6'b111111;
mem[38] = 6'b111111;
mem[39] = 6'b111111;
mem[40] = 6'b111111;
mem[41] = 6'b111111;
mem[42] = 6'b111111;
mem[43] = 6'b111111;
mem[44] = 6'b111111;
mem[45] = 6'b111111;
mem[46] = 6'b111111;
mem[47] = 6'b111111;
mem[48] = 6'b111111;
mem[49] = 6'b111111;
mem[50] = 6'b111111;
mem[51] = 6'b111111;
mem[52] = 6'b111111;
mem[53] = 6'b111111;
mem[54] = 6'b111111;
mem[55] = 6'b111111;
mem[56] = 6'b111111;
mem[57] = 6'b111111;
mem[58] = 6'b111111;
mem[59] = 6'b111111;
mem[60] = 6'b111111;
mem[61] = 6'b111111;
mem[62] = 6'b111111;
mem[63] = 6'b111111;
mem[64] = 6'b111111;
mem[65] = 6'b111111;
mem[66] = 6'b111111;
mem[67] = 6'b111111;
mem[68] = 6'b111111;
mem[69] = 6'b111111;
mem[70] = 6'b111111;
mem[71] = 6'b111111;
mem[72] = 6'b111111;
mem[73] = 6'b111111;
mem[74] = 6'b111111;
mem[75] = 6'b111111;
mem[76] = 6'b111111;
mem[77] = 6'b111111;
mem[78] = 6'b111111;
mem[79] = 6'b111111;
mem[80] = 6'b111111;
mem[81] = 6'b111111;
mem[82] = 6'b111111;
mem[83] = 6'b111111;
mem[84] = 6'b111111;
mem[85] = 6'b111111;
mem[86] = 6'b111111;
mem[87] = 6'b111111;
mem[88] = 6'b111111;
mem[89] = 6'b111111;
mem[90] = 6'b111111;
mem[91] = 6'b111111;
mem[92] = 6'b111111;
mem[93] = 6'b111111;
mem[94] = 6'b111111;
mem[95] = 6'b111111;
mem[96] = 6'b111111;
mem[97] = 6'b111111;
mem[98] = 6'b111111;
mem[99] = 6'b111111;
mem[100] = 6'b111111;
mem[101] = 6'b111111;
mem[102] = 6'b111111;
mem[103] = 6'b111111;
mem[104] = 6'b111111;
mem[105] = 6'b111111;
mem[106] = 6'b111111;
mem[107] = 6'b111111;
mem[108] = 6'b111111;
mem[109] = 6'b111111;
mem[110] = 6'b111111;
mem[111] = 6'b111111;
mem[112] = 6'b111111;
mem[113] = 6'b111111;
mem[114] = 6'b111111;
mem[115] = 6'b111111;
mem[116] = 6'b111111;
mem[117] = 6'b111111;
mem[118] = 6'b111111;
mem[119] = 6'b111111;
mem[120] = 6'b111111;
mem[121] = 6'b111111;
mem[122] = 6'b111111;
mem[123] = 6'b111111;
mem[124] = 6'b111111;
mem[125] = 6'b111111;
mem[126] = 6'b111111;
mem[127] = 6'b111111;
mem[128] = 6'b111111;
mem[129] = 6'b111111;
mem[130] = 6'b111111;
mem[131] = 6'b111111;
mem[132] = 6'b111111;
mem[133] = 6'b111111;
mem[134] = 6'b111111;
mem[135] = 6'b111111;
mem[136] = 6'b111111;
mem[137] = 6'b111111;
mem[138] = 6'b111111;
mem[139] = 6'b111111;
mem[140] = 6'b111111;
mem[141] = 6'b111111;
mem[142] = 6'b111111;
mem[143] = 6'b111111;
mem[144] = 6'b111111;
mem[145] = 6'b111111;
mem[146] = 6'b111111;
mem[147] = 6'b111111;
mem[148] = 6'b111111;
mem[149] = 6'b111111;
mem[150] = 6'b111111;
mem[151] = 6'b111111;
mem[152] = 6'b111111;
mem[153] = 6'b111111;
mem[154] = 6'b111111;
mem[155] = 6'b111111;
mem[156] = 6'b111111;
mem[157] = 6'b111111;
mem[158] = 6'b111111;
mem[159] = 6'b111111;
mem[160] = 6'b111111;
mem[161] = 6'b111111;
mem[162] = 6'b111111;
mem[163] = 6'b111111;
mem[164] = 6'b111111;
mem[165] = 6'b111111;
mem[166] = 6'b111111;
mem[167] = 6'b111111;
mem[168] = 6'b111111;
mem[169] = 6'b111111;
mem[170] = 6'b111111;
mem[171] = 6'b111111;
mem[172] = 6'b111111;
mem[173] = 6'b111111;
mem[174] = 6'b111111;
mem[175] = 6'b111111;
mem[176] = 6'b111111;
mem[177] = 6'b111111;
mem[178] = 6'b111111;
mem[179] = 6'b111111;
mem[180] = 6'b111111;
mem[181] = 6'b111111;
mem[182] = 6'b111111;
mem[183] = 6'b111111;
mem[184] = 6'b111111;
mem[185] = 6'b111111;
mem[186] = 6'b111111;
mem[187] = 6'b111111;
mem[188] = 6'b111111;
mem[189] = 6'b111111;
mem[190] = 6'b111111;
mem[191] = 6'b111111;
mem[192] = 6'b111111;
mem[193] = 6'b111111;
mem[194] = 6'b111111;
mem[195] = 6'b111111;
mem[196] = 6'b111111;
mem[197] = 6'b111111;
mem[198] = 6'b111111;
mem[199] = 6'b111111;
mem[200] = 6'b111111;
mem[201] = 6'b111111;
mem[202] = 6'b111111;
mem[203] = 6'b111111;
mem[204] = 6'b111111;
mem[205] = 6'b111111;
mem[206] = 6'b111111;
mem[207] = 6'b111111;
mem[208] = 6'b111111;
mem[209] = 6'b111111;
mem[210] = 6'b111111;
mem[211] = 6'b111111;
mem[212] = 6'b111111;
mem[213] = 6'b111111;
mem[214] = 6'b111111;
mem[215] = 6'b111111;
mem[216] = 6'b111111;
mem[217] = 6'b111111;
mem[218] = 6'b111111;
mem[219] = 6'b111111;
mem[220] = 6'b111111;
mem[221] = 6'b111111;
mem[222] = 6'b111111;
mem[223] = 6'b111111;
mem[224] = 6'b111111;
mem[225] = 6'b111111;
mem[226] = 6'b111111;
mem[227] = 6'b111111;
mem[228] = 6'b111111;
mem[229] = 6'b111111;
mem[230] = 6'b111111;
mem[231] = 6'b111111;
mem[232] = 6'b111111;
mem[233] = 6'b111111;
mem[234] = 6'b111111;
mem[235] = 6'b111111;
mem[236] = 6'b111111;
mem[237] = 6'b111111;
mem[238] = 6'b111111;
mem[239] = 6'b111111;
mem[240] = 6'b111111;
mem[241] = 6'b111111;
mem[242] = 6'b111111;
mem[243] = 6'b111111;
mem[244] = 6'b111111;
mem[245] = 6'b111111;
mem[246] = 6'b111111;
mem[247] = 6'b111111;
mem[248] = 6'b111111;
mem[249] = 6'b111111;
mem[250] = 6'b111111;
mem[251] = 6'b111111;
mem[252] = 6'b111111;
mem[253] = 6'b111111;
mem[254] = 6'b111111;
mem[255] = 6'b111111;
mem[256] = 6'b111111;
mem[257] = 6'b111111;
mem[258] = 6'b111111;
mem[259] = 6'b111111;
mem[260] = 6'b111111;
mem[261] = 6'b111111;
mem[262] = 6'b111111;
mem[263] = 6'b111111;
mem[264] = 6'b111111;
mem[265] = 6'b111111;
mem[266] = 6'b111111;
mem[267] = 6'b111111;
mem[268] = 6'b111111;
mem[269] = 6'b111111;
mem[270] = 6'b111111;
mem[271] = 6'b111111;
mem[272] = 6'b111111;
mem[273] = 6'b111111;
mem[274] = 6'b111111;
mem[275] = 6'b111111;
mem[276] = 6'b111111;
mem[277] = 6'b111111;
mem[278] = 6'b111111;
mem[279] = 6'b111111;
mem[280] = 6'b111111;
mem[281] = 6'b111111;
mem[282] = 6'b111111;
mem[283] = 6'b111111;
mem[284] = 6'b111111;
mem[285] = 6'b111111;
mem[286] = 6'b111111;
mem[287] = 6'b111111;
mem[288] = 6'b111111;
mem[289] = 6'b111111;
mem[290] = 6'b111111;
mem[291] = 6'b111111;
mem[292] = 6'b111111;
mem[293] = 6'b111111;
mem[294] = 6'b111111;
mem[295] = 6'b111111;
mem[296] = 6'b111111;
mem[297] = 6'b111111;
mem[298] = 6'b111111;
mem[299] = 6'b111111;
mem[300] = 6'b111111;
mem[301] = 6'b111111;
mem[302] = 6'b111111;
mem[303] = 6'b111111;
mem[304] = 6'b111111;
mem[305] = 6'b111111;
mem[306] = 6'b111111;
mem[307] = 6'b111111;
mem[308] = 6'b111111;
mem[309] = 6'b111111;
mem[310] = 6'b111111;
mem[311] = 6'b111111;
mem[312] = 6'b111111;
mem[313] = 6'b111111;
mem[314] = 6'b111111;
mem[315] = 6'b111111;
mem[316] = 6'b111111;
mem[317] = 6'b111111;
mem[318] = 6'b111111;
mem[319] = 6'b111111;
mem[320] = 6'b111111;
mem[321] = 6'b111111;
mem[322] = 6'b111111;
mem[323] = 6'b111111;
mem[324] = 6'b111111;
mem[325] = 6'b111111;
mem[326] = 6'b111111;
mem[327] = 6'b111111;
mem[328] = 6'b111111;
mem[329] = 6'b111111;
mem[330] = 6'b111111;
mem[331] = 6'b111111;
mem[332] = 6'b111111;
mem[333] = 6'b111111;
mem[334] = 6'b111111;
mem[335] = 6'b111111;
mem[336] = 6'b111111;
mem[337] = 6'b111111;
mem[338] = 6'b111111;
mem[339] = 6'b111111;
mem[340] = 6'b111111;
mem[341] = 6'b111111;
mem[342] = 6'b111111;
mem[343] = 6'b111111;
mem[344] = 6'b111111;
mem[345] = 6'b111111;
mem[346] = 6'b111111;
mem[347] = 6'b111111;
mem[348] = 6'b111111;
mem[349] = 6'b111111;
mem[350] = 6'b111111;
mem[351] = 6'b111111;
mem[352] = 6'b111111;
mem[353] = 6'b111111;
mem[354] = 6'b111111;
mem[355] = 6'b111111;
mem[356] = 6'b111111;
mem[357] = 6'b111111;
mem[358] = 6'b111111;
mem[359] = 6'b111111;
mem[360] = 6'b111111;
mem[361] = 6'b111111;
mem[362] = 6'b111111;
mem[363] = 6'b111111;
mem[364] = 6'b111111;
mem[365] = 6'b111111;
mem[366] = 6'b111111;
mem[367] = 6'b111111;
mem[368] = 6'b111111;
mem[369] = 6'b111111;
mem[370] = 6'b111111;
mem[371] = 6'b111111;
mem[372] = 6'b111111;
mem[373] = 6'b111111;
mem[374] = 6'b111111;
mem[375] = 6'b111111;
mem[376] = 6'b111111;
mem[377] = 6'b111111;
mem[378] = 6'b111111;
mem[379] = 6'b111111;
mem[380] = 6'b111111;
mem[381] = 6'b111111;
mem[382] = 6'b111111;
mem[383] = 6'b111111;
mem[384] = 6'b111111;
mem[385] = 6'b111111;
mem[386] = 6'b111111;
mem[387] = 6'b111111;
mem[388] = 6'b111111;
mem[389] = 6'b111111;
mem[390] = 6'b111111;
mem[391] = 6'b111111;
mem[392] = 6'b111111;
mem[393] = 6'b111111;
mem[394] = 6'b111111;
mem[395] = 6'b111111;
mem[396] = 6'b111111;
mem[397] = 6'b111111;
mem[398] = 6'b111111;
mem[399] = 6'b111111;
mem[400] = 6'b111111;
mem[401] = 6'b111111;
mem[402] = 6'b111111;
mem[403] = 6'b111111;
mem[404] = 6'b111111;
mem[405] = 6'b111111;
mem[406] = 6'b111111;
mem[407] = 6'b111111;
mem[408] = 6'b111111;
mem[409] = 6'b111111;
mem[410] = 6'b111111;
mem[411] = 6'b111111;
mem[412] = 6'b111111;
mem[413] = 6'b111111;
mem[414] = 6'b111111;
mem[415] = 6'b111111;
mem[416] = 6'b111111;
mem[417] = 6'b111111;
mem[418] = 6'b111111;
mem[419] = 6'b111111;
mem[420] = 6'b111111;
mem[421] = 6'b111111;
mem[422] = 6'b111111;
mem[423] = 6'b111111;
mem[424] = 6'b111111;
mem[425] = 6'b111111;
mem[426] = 6'b111111;
mem[427] = 6'b111111;
mem[428] = 6'b111111;
mem[429] = 6'b111111;
mem[430] = 6'b111111;
mem[431] = 6'b111111;
mem[432] = 6'b111111;
mem[433] = 6'b111111;
mem[434] = 6'b111111;
mem[435] = 6'b111111;
mem[436] = 6'b111111;
mem[437] = 6'b111111;
mem[438] = 6'b111111;
mem[439] = 6'b111111;
mem[440] = 6'b111111;
mem[441] = 6'b111111;
mem[442] = 6'b111111;
mem[443] = 6'b111111;
mem[444] = 6'b111111;
mem[445] = 6'b111111;
mem[446] = 6'b111111;
mem[447] = 6'b111111;
mem[448] = 6'b111111;
mem[449] = 6'b111111;
mem[450] = 6'b111111;
mem[451] = 6'b111111;
mem[452] = 6'b111111;
mem[453] = 6'b111111;
mem[454] = 6'b111111;
mem[455] = 6'b111111;
mem[456] = 6'b111111;
mem[457] = 6'b111111;
mem[458] = 6'b111111;
mem[459] = 6'b111111;
mem[460] = 6'b111111;
mem[461] = 6'b111111;
mem[462] = 6'b111111;
mem[463] = 6'b111111;
mem[464] = 6'b111111;
mem[465] = 6'b111111;
mem[466] = 6'b111111;
mem[467] = 6'b111111;
mem[468] = 6'b111111;
mem[469] = 6'b111111;
mem[470] = 6'b111111;
mem[471] = 6'b111111;
mem[472] = 6'b111111;
mem[473] = 6'b111111;
mem[474] = 6'b111111;
mem[475] = 6'b111111;
mem[476] = 6'b111111;
mem[477] = 6'b111111;
mem[478] = 6'b111111;
mem[479] = 6'b111111;
mem[480] = 6'b111111;
mem[481] = 6'b111111;
mem[482] = 6'b111111;
mem[483] = 6'b111111;
mem[484] = 6'b111111;
mem[485] = 6'b111111;
mem[486] = 6'b111111;
mem[487] = 6'b111111;
mem[488] = 6'b111111;
mem[489] = 6'b111111;
mem[490] = 6'b111111;
mem[491] = 6'b111111;
mem[492] = 6'b111111;
mem[493] = 6'b111111;
mem[494] = 6'b111111;
mem[495] = 6'b111111;
mem[496] = 6'b111111;
mem[497] = 6'b111111;
mem[498] = 6'b111111;
mem[499] = 6'b111111;
mem[500] = 6'b111111;
mem[501] = 6'b111111;
mem[502] = 6'b111111;
mem[503] = 6'b111111;
mem[504] = 6'b111111;
mem[505] = 6'b111111;
mem[506] = 6'b111111;
mem[507] = 6'b111111;
mem[508] = 6'b111111;
mem[509] = 6'b111111;
mem[510] = 6'b111111;
mem[511] = 6'b111111;
mem[512] = 6'b111111;
mem[513] = 6'b111111;
mem[514] = 6'b111111;
mem[515] = 6'b111111;
mem[516] = 6'b111111;
mem[517] = 6'b111111;
mem[518] = 6'b111111;
mem[519] = 6'b111111;
mem[520] = 6'b111111;
mem[521] = 6'b111111;
mem[522] = 6'b111111;
mem[523] = 6'b111111;
mem[524] = 6'b111111;
mem[525] = 6'b111111;
mem[526] = 6'b111111;
mem[527] = 6'b111111;
mem[528] = 6'b111111;
mem[529] = 6'b111111;
mem[530] = 6'b111111;
mem[531] = 6'b111111;
mem[532] = 6'b111111;
mem[533] = 6'b111111;
mem[534] = 6'b111111;
mem[535] = 6'b111111;
mem[536] = 6'b111111;
mem[537] = 6'b111111;
mem[538] = 6'b111111;
mem[539] = 6'b111111;
mem[540] = 6'b111111;
mem[541] = 6'b111111;
mem[542] = 6'b111111;
mem[543] = 6'b111111;
mem[544] = 6'b111111;
mem[545] = 6'b101010;
mem[546] = 6'b011010;
mem[547] = 6'b111111;
mem[548] = 6'b111111;
mem[549] = 6'b111111;
mem[550] = 6'b111111;
mem[551] = 6'b111111;
mem[552] = 6'b111111;
mem[553] = 6'b111111;
mem[554] = 6'b111111;
mem[555] = 6'b111111;
mem[556] = 6'b111111;
mem[557] = 6'b111111;
mem[558] = 6'b111111;
mem[559] = 6'b111111;
mem[560] = 6'b111111;
mem[561] = 6'b111111;
mem[562] = 6'b111111;
mem[563] = 6'b111111;
mem[564] = 6'b111111;
mem[565] = 6'b111111;
mem[566] = 6'b111111;
mem[567] = 6'b111111;
mem[568] = 6'b111111;
mem[569] = 6'b111111;
mem[570] = 6'b111111;
mem[571] = 6'b111111;
mem[572] = 6'b111111;
mem[573] = 6'b111111;
mem[574] = 6'b111111;
mem[575] = 6'b111111;
mem[576] = 6'b111111;
mem[577] = 6'b111111;
mem[578] = 6'b111111;
mem[579] = 6'b111111;
mem[580] = 6'b111111;
mem[581] = 6'b111111;
mem[582] = 6'b111111;
mem[583] = 6'b111111;
mem[584] = 6'b111111;
mem[585] = 6'b111111;
mem[586] = 6'b111111;
mem[587] = 6'b111111;
mem[588] = 6'b111111;
mem[589] = 6'b111111;
mem[590] = 6'b111111;
mem[591] = 6'b111111;
mem[592] = 6'b111111;
mem[593] = 6'b111111;
mem[594] = 6'b111111;
mem[595] = 6'b111111;
mem[596] = 6'b111111;
mem[597] = 6'b111111;
mem[598] = 6'b111111;
mem[599] = 6'b111111;
mem[600] = 6'b111111;
mem[601] = 6'b101010;
mem[602] = 6'b001001;
mem[603] = 6'b111111;
mem[604] = 6'b000101;
mem[605] = 6'b111111;
mem[606] = 6'b000101;
mem[607] = 6'b000101;
mem[608] = 6'b001001;
mem[609] = 6'b000101;
mem[610] = 6'b000101;
mem[611] = 6'b101010;
mem[612] = 6'b000101;
mem[613] = 6'b011010;
mem[614] = 6'b001001;
mem[615] = 6'b111111;
mem[616] = 6'b111111;
mem[617] = 6'b111111;
mem[618] = 6'b111111;
mem[619] = 6'b111111;
mem[620] = 6'b111111;
mem[621] = 6'b111111;
mem[622] = 6'b111111;
mem[623] = 6'b111111;
mem[624] = 6'b111111;
mem[625] = 6'b111111;
mem[626] = 6'b111111;
mem[627] = 6'b111111;
mem[628] = 6'b111111;
mem[629] = 6'b111111;
mem[630] = 6'b111111;
mem[631] = 6'b111111;
mem[632] = 6'b111111;
mem[633] = 6'b111111;
mem[634] = 6'b111111;
mem[635] = 6'b111111;
mem[636] = 6'b111111;
mem[637] = 6'b111111;
mem[638] = 6'b111111;
mem[639] = 6'b111111;
mem[640] = 6'b111111;
mem[641] = 6'b111111;
mem[642] = 6'b111111;
mem[643] = 6'b111111;
mem[644] = 6'b111111;
mem[645] = 6'b111111;
mem[646] = 6'b111111;
mem[647] = 6'b111111;
mem[648] = 6'b111111;
mem[649] = 6'b111111;
mem[650] = 6'b111111;
mem[651] = 6'b111111;
mem[652] = 6'b111111;
mem[653] = 6'b111111;
mem[654] = 6'b111111;
mem[655] = 6'b111111;
mem[656] = 6'b111111;
mem[657] = 6'b111111;
mem[658] = 6'b111111;
mem[659] = 6'b111111;
mem[660] = 6'b111111;
mem[661] = 6'b111111;
mem[662] = 6'b111111;
mem[663] = 6'b011010;
mem[664] = 6'b011010;
mem[665] = 6'b000101;
mem[666] = 6'b000101;
mem[667] = 6'b011010;
mem[668] = 6'b000101;
mem[669] = 6'b011010;
mem[670] = 6'b000101;
mem[671] = 6'b011010;
mem[672] = 6'b111111;
mem[673] = 6'b000101;
mem[674] = 6'b000101;
mem[675] = 6'b011010;
mem[676] = 6'b001001;
mem[677] = 6'b000101;
mem[678] = 6'b101010;
mem[679] = 6'b000101;
mem[680] = 6'b000101;
mem[681] = 6'b111111;
mem[682] = 6'b111111;
mem[683] = 6'b111111;
mem[684] = 6'b111111;
mem[685] = 6'b111111;
mem[686] = 6'b111111;
mem[687] = 6'b111111;
mem[688] = 6'b111111;
mem[689] = 6'b111111;
mem[690] = 6'b111111;
mem[691] = 6'b111111;
mem[692] = 6'b111111;
mem[693] = 6'b111111;
mem[694] = 6'b111111;
mem[695] = 6'b111111;
mem[696] = 6'b111111;
mem[697] = 6'b111111;
mem[698] = 6'b111111;
mem[699] = 6'b111111;
mem[700] = 6'b111111;
mem[701] = 6'b111111;
mem[702] = 6'b111111;
mem[703] = 6'b111111;
mem[704] = 6'b111111;
mem[705] = 6'b111111;
mem[706] = 6'b111111;
mem[707] = 6'b111111;
mem[708] = 6'b111111;
mem[709] = 6'b111111;
mem[710] = 6'b111111;
mem[711] = 6'b111111;
mem[712] = 6'b111111;
mem[713] = 6'b111111;
mem[714] = 6'b111111;
mem[715] = 6'b111111;
mem[716] = 6'b111111;
mem[717] = 6'b111111;
mem[718] = 6'b111111;
mem[719] = 6'b111111;
mem[720] = 6'b111111;
mem[721] = 6'b111111;
mem[722] = 6'b111111;
mem[723] = 6'b111111;
mem[724] = 6'b111111;
mem[725] = 6'b000101;
mem[726] = 6'b101010;
mem[727] = 6'b101010;
mem[728] = 6'b101010;
mem[729] = 6'b000101;
mem[730] = 6'b000101;
mem[731] = 6'b011010;
mem[732] = 6'b000101;
mem[733] = 6'b001001;
mem[734] = 6'b101010;
mem[735] = 6'b101010;
mem[736] = 6'b000101;
mem[737] = 6'b111111;
mem[738] = 6'b111111;
mem[739] = 6'b000101;
mem[740] = 6'b000101;
mem[741] = 6'b000101;
mem[742] = 6'b101010;
mem[743] = 6'b000101;
mem[744] = 6'b000101;
mem[745] = 6'b111111;
mem[746] = 6'b000101;
mem[747] = 6'b111111;
mem[748] = 6'b111111;
mem[749] = 6'b111111;
mem[750] = 6'b111111;
mem[751] = 6'b111111;
mem[752] = 6'b111111;
mem[753] = 6'b111111;
mem[754] = 6'b111111;
mem[755] = 6'b111111;
mem[756] = 6'b111111;
mem[757] = 6'b111111;
mem[758] = 6'b111111;
mem[759] = 6'b111111;
mem[760] = 6'b111111;
mem[761] = 6'b111111;
mem[762] = 6'b111111;
mem[763] = 6'b111111;
mem[764] = 6'b111111;
mem[765] = 6'b111111;
mem[766] = 6'b111111;
mem[767] = 6'b111111;
mem[768] = 6'b111111;
mem[769] = 6'b111111;
mem[770] = 6'b111111;
mem[771] = 6'b111111;
mem[772] = 6'b111111;
mem[773] = 6'b111111;
mem[774] = 6'b111111;
mem[775] = 6'b111111;
mem[776] = 6'b111111;
mem[777] = 6'b111111;
mem[778] = 6'b111111;
mem[779] = 6'b111111;
mem[780] = 6'b111111;
mem[781] = 6'b111111;
mem[782] = 6'b111111;
mem[783] = 6'b111111;
mem[784] = 6'b111111;
mem[785] = 6'b111111;
mem[786] = 6'b111111;
mem[787] = 6'b011001;
mem[788] = 6'b000101;
mem[789] = 6'b101010;
mem[790] = 6'b000101;
mem[791] = 6'b000101;
mem[792] = 6'b001001;
mem[793] = 6'b011010;
mem[794] = 6'b000101;
mem[795] = 6'b000101;
mem[796] = 6'b000101;
mem[797] = 6'b000101;
mem[798] = 6'b000101;
mem[799] = 6'b000101;
mem[800] = 6'b000101;
mem[801] = 6'b000101;
mem[802] = 6'b000101;
mem[803] = 6'b111111;
mem[804] = 6'b000101;
mem[805] = 6'b001001;
mem[806] = 6'b011010;
mem[807] = 6'b101010;
mem[808] = 6'b101010;
mem[809] = 6'b000101;
mem[810] = 6'b001001;
mem[811] = 6'b011001;
mem[812] = 6'b000101;
mem[813] = 6'b101010;
mem[814] = 6'b111111;
mem[815] = 6'b111111;
mem[816] = 6'b111111;
mem[817] = 6'b111111;
mem[818] = 6'b111111;
mem[819] = 6'b111111;
mem[820] = 6'b111111;
mem[821] = 6'b111111;
mem[822] = 6'b111111;
mem[823] = 6'b111111;
mem[824] = 6'b111111;
mem[825] = 6'b111111;
mem[826] = 6'b111111;
mem[827] = 6'b111111;
mem[828] = 6'b111111;
mem[829] = 6'b111111;
mem[830] = 6'b111111;
mem[831] = 6'b111111;
mem[832] = 6'b111111;
mem[833] = 6'b111111;
mem[834] = 6'b111111;
mem[835] = 6'b111111;
mem[836] = 6'b111111;
mem[837] = 6'b111111;
mem[838] = 6'b111111;
mem[839] = 6'b111111;
mem[840] = 6'b111111;
mem[841] = 6'b111111;
mem[842] = 6'b111111;
mem[843] = 6'b111111;
mem[844] = 6'b111111;
mem[845] = 6'b111111;
mem[846] = 6'b111111;
mem[847] = 6'b111111;
mem[848] = 6'b111111;
mem[849] = 6'b111111;
mem[850] = 6'b000101;
mem[851] = 6'b000101;
mem[852] = 6'b000101;
mem[853] = 6'b000101;
mem[854] = 6'b101010;
mem[855] = 6'b000101;
mem[856] = 6'b011010;
mem[857] = 6'b001001;
mem[858] = 6'b000101;
mem[859] = 6'b111111;
mem[860] = 6'b001001;
mem[861] = 6'b111111;
mem[862] = 6'b101010;
mem[863] = 6'b101010;
mem[864] = 6'b001001;
mem[865] = 6'b101010;
mem[866] = 6'b101010;
mem[867] = 6'b101010;
mem[868] = 6'b000101;
mem[869] = 6'b000101;
mem[870] = 6'b101010;
mem[871] = 6'b000101;
mem[872] = 6'b011010;
mem[873] = 6'b111111;
mem[874] = 6'b011010;
mem[875] = 6'b000101;
mem[876] = 6'b000101;
mem[877] = 6'b000101;
mem[878] = 6'b111111;
mem[879] = 6'b111111;
mem[880] = 6'b111111;
mem[881] = 6'b111111;
mem[882] = 6'b111111;
mem[883] = 6'b111111;
mem[884] = 6'b111111;
mem[885] = 6'b111111;
mem[886] = 6'b111111;
mem[887] = 6'b111111;
mem[888] = 6'b111111;
mem[889] = 6'b111111;
mem[890] = 6'b111111;
mem[891] = 6'b111111;
mem[892] = 6'b111111;
mem[893] = 6'b111111;
mem[894] = 6'b111111;
mem[895] = 6'b111111;
mem[896] = 6'b111111;
mem[897] = 6'b111111;
mem[898] = 6'b111111;
mem[899] = 6'b111111;
mem[900] = 6'b111111;
mem[901] = 6'b111111;
mem[902] = 6'b111111;
mem[903] = 6'b111111;
mem[904] = 6'b111111;
mem[905] = 6'b111111;
mem[906] = 6'b111111;
mem[907] = 6'b111111;
mem[908] = 6'b111111;
mem[909] = 6'b111111;
mem[910] = 6'b111111;
mem[911] = 6'b111111;
mem[912] = 6'b111111;
mem[913] = 6'b111111;
mem[914] = 6'b001001;
mem[915] = 6'b101010;
mem[916] = 6'b001001;
mem[917] = 6'b101010;
mem[918] = 6'b101010;
mem[919] = 6'b000101;
mem[920] = 6'b001001;
mem[921] = 6'b101010;
mem[922] = 6'b101010;
mem[923] = 6'b000101;
mem[924] = 6'b111111;
mem[925] = 6'b000101;
mem[926] = 6'b011001;
mem[927] = 6'b000101;
mem[928] = 6'b000101;
mem[929] = 6'b101010;
mem[930] = 6'b000101;
mem[931] = 6'b001001;
mem[932] = 6'b000101;
mem[933] = 6'b000101;
mem[934] = 6'b111111;
mem[935] = 6'b101010;
mem[936] = 6'b101010;
mem[937] = 6'b000101;
mem[938] = 6'b111111;
mem[939] = 6'b101010;
mem[940] = 6'b000101;
mem[941] = 6'b101010;
mem[942] = 6'b000101;
mem[943] = 6'b111111;
mem[944] = 6'b111111;
mem[945] = 6'b111111;
mem[946] = 6'b111111;
mem[947] = 6'b111111;
mem[948] = 6'b111111;
mem[949] = 6'b111111;
mem[950] = 6'b111111;
mem[951] = 6'b111111;
mem[952] = 6'b111111;
mem[953] = 6'b111111;
mem[954] = 6'b111111;
mem[955] = 6'b111111;
mem[956] = 6'b111111;
mem[957] = 6'b111111;
mem[958] = 6'b111111;
mem[959] = 6'b111111;
mem[960] = 6'b111111;
mem[961] = 6'b111111;
mem[962] = 6'b111111;
mem[963] = 6'b111111;
mem[964] = 6'b111111;
mem[965] = 6'b111111;
mem[966] = 6'b111111;
mem[967] = 6'b111111;
mem[968] = 6'b111111;
mem[969] = 6'b111111;
mem[970] = 6'b111111;
mem[971] = 6'b111111;
mem[972] = 6'b111111;
mem[973] = 6'b111111;
mem[974] = 6'b111111;
mem[975] = 6'b111111;
mem[976] = 6'b011010;
mem[977] = 6'b001001;
mem[978] = 6'b000101;
mem[979] = 6'b000101;
mem[980] = 6'b101010;
mem[981] = 6'b000101;
mem[982] = 6'b011010;
mem[983] = 6'b111111;
mem[984] = 6'b000101;
mem[985] = 6'b000101;
mem[986] = 6'b101010;
mem[987] = 6'b000101;
mem[988] = 6'b101010;
mem[989] = 6'b011010;
mem[990] = 6'b111111;
mem[991] = 6'b000101;
mem[992] = 6'b000101;
mem[993] = 6'b111111;
mem[994] = 6'b011010;
mem[995] = 6'b111111;
mem[996] = 6'b000101;
mem[997] = 6'b001001;
mem[998] = 6'b000101;
mem[999] = 6'b101010;
mem[1000] = 6'b000101;
mem[1001] = 6'b000101;
mem[1002] = 6'b000101;
mem[1003] = 6'b000101;
mem[1004] = 6'b011010;
mem[1005] = 6'b101010;
mem[1006] = 6'b101010;
mem[1007] = 6'b101010;
mem[1008] = 6'b111111;
mem[1009] = 6'b111111;
mem[1010] = 6'b111111;
mem[1011] = 6'b111111;
mem[1012] = 6'b111111;
mem[1013] = 6'b111111;
mem[1014] = 6'b111111;
mem[1015] = 6'b111111;
mem[1016] = 6'b111111;
mem[1017] = 6'b111111;
mem[1018] = 6'b111111;
mem[1019] = 6'b111111;
mem[1020] = 6'b111111;
mem[1021] = 6'b111111;
mem[1022] = 6'b111111;
mem[1023] = 6'b111111;
mem[1024] = 6'b111111;
mem[1025] = 6'b111111;
mem[1026] = 6'b111111;
mem[1027] = 6'b111111;
mem[1028] = 6'b111111;
mem[1029] = 6'b111111;
mem[1030] = 6'b111111;
mem[1031] = 6'b111111;
mem[1032] = 6'b111111;
mem[1033] = 6'b111111;
mem[1034] = 6'b111111;
mem[1035] = 6'b111111;
mem[1036] = 6'b111111;
mem[1037] = 6'b111111;
mem[1038] = 6'b111111;
mem[1039] = 6'b000101;
mem[1040] = 6'b000101;
mem[1041] = 6'b101010;
mem[1042] = 6'b000101;
mem[1043] = 6'b000101;
mem[1044] = 6'b101010;
mem[1045] = 6'b011010;
mem[1046] = 6'b101111;
mem[1047] = 6'b111111;
mem[1048] = 6'b000101;
mem[1049] = 6'b000101;
mem[1050] = 6'b000101;
mem[1051] = 6'b011010;
mem[1052] = 6'b000101;
mem[1053] = 6'b111111;
mem[1054] = 6'b001001;
mem[1055] = 6'b000101;
mem[1056] = 6'b000101;
mem[1057] = 6'b111111;
mem[1058] = 6'b000101;
mem[1059] = 6'b011010;
mem[1060] = 6'b011010;
mem[1061] = 6'b101010;
mem[1062] = 6'b011010;
mem[1063] = 6'b111111;
mem[1064] = 6'b011010;
mem[1065] = 6'b000101;
mem[1066] = 6'b111111;
mem[1067] = 6'b001001;
mem[1068] = 6'b111111;
mem[1069] = 6'b000101;
mem[1070] = 6'b000101;
mem[1071] = 6'b001001;
mem[1072] = 6'b000101;
mem[1073] = 6'b111111;
mem[1074] = 6'b111111;
mem[1075] = 6'b111111;
mem[1076] = 6'b111111;
mem[1077] = 6'b111111;
mem[1078] = 6'b111111;
mem[1079] = 6'b111111;
mem[1080] = 6'b111111;
mem[1081] = 6'b111111;
mem[1082] = 6'b111111;
mem[1083] = 6'b111111;
mem[1084] = 6'b111111;
mem[1085] = 6'b111111;
mem[1086] = 6'b111111;
mem[1087] = 6'b111111;
mem[1088] = 6'b111111;
mem[1089] = 6'b111111;
mem[1090] = 6'b111111;
mem[1091] = 6'b111111;
mem[1092] = 6'b111111;
mem[1093] = 6'b111111;
mem[1094] = 6'b111111;
mem[1095] = 6'b111111;
mem[1096] = 6'b111111;
mem[1097] = 6'b111111;
mem[1098] = 6'b111111;
mem[1099] = 6'b111111;
mem[1100] = 6'b111111;
mem[1101] = 6'b111111;
mem[1102] = 6'b000101;
mem[1103] = 6'b101010;
mem[1104] = 6'b011010;
mem[1105] = 6'b000101;
mem[1106] = 6'b000101;
mem[1107] = 6'b011010;
mem[1108] = 6'b000101;
mem[1109] = 6'b000101;
mem[1110] = 6'b000101;
mem[1111] = 6'b101010;
mem[1112] = 6'b111111;
mem[1113] = 6'b011010;
mem[1114] = 6'b011010;
mem[1115] = 6'b000101;
mem[1116] = 6'b000101;
mem[1117] = 6'b000101;
mem[1118] = 6'b000101;
mem[1119] = 6'b011010;
mem[1120] = 6'b111111;
mem[1121] = 6'b011010;
mem[1122] = 6'b000101;
mem[1123] = 6'b101010;
mem[1124] = 6'b000101;
mem[1125] = 6'b000101;
mem[1126] = 6'b101010;
mem[1127] = 6'b000101;
mem[1128] = 6'b111111;
mem[1129] = 6'b000101;
mem[1130] = 6'b000101;
mem[1131] = 6'b000101;
mem[1132] = 6'b101010;
mem[1133] = 6'b000101;
mem[1134] = 6'b000101;
mem[1135] = 6'b111111;
mem[1136] = 6'b101010;
mem[1137] = 6'b000101;
mem[1138] = 6'b111111;
mem[1139] = 6'b111111;
mem[1140] = 6'b111111;
mem[1141] = 6'b111111;
mem[1142] = 6'b111111;
mem[1143] = 6'b111111;
mem[1144] = 6'b111111;
mem[1145] = 6'b111111;
mem[1146] = 6'b111111;
mem[1147] = 6'b111111;
mem[1148] = 6'b111111;
mem[1149] = 6'b111111;
mem[1150] = 6'b111111;
mem[1151] = 6'b111111;
mem[1152] = 6'b111111;
mem[1153] = 6'b111111;
mem[1154] = 6'b111111;
mem[1155] = 6'b111111;
mem[1156] = 6'b111111;
mem[1157] = 6'b111111;
mem[1158] = 6'b111111;
mem[1159] = 6'b111111;
mem[1160] = 6'b111111;
mem[1161] = 6'b111111;
mem[1162] = 6'b111111;
mem[1163] = 6'b111111;
mem[1164] = 6'b111111;
mem[1165] = 6'b101010;
mem[1166] = 6'b101010;
mem[1167] = 6'b000101;
mem[1168] = 6'b000101;
mem[1169] = 6'b000101;
mem[1170] = 6'b000101;
mem[1171] = 6'b011010;
mem[1172] = 6'b000101;
mem[1173] = 6'b000101;
mem[1174] = 6'b011010;
mem[1175] = 6'b001001;
mem[1176] = 6'b000101;
mem[1177] = 6'b001001;
mem[1178] = 6'b011001;
mem[1179] = 6'b101010;
mem[1180] = 6'b000101;
mem[1181] = 6'b001001;
mem[1182] = 6'b000101;
mem[1183] = 6'b011010;
mem[1184] = 6'b000101;
mem[1185] = 6'b000101;
mem[1186] = 6'b001001;
mem[1187] = 6'b111111;
mem[1188] = 6'b000101;
mem[1189] = 6'b000101;
mem[1190] = 6'b111111;
mem[1191] = 6'b101010;
mem[1192] = 6'b100101;
mem[1193] = 6'b111111;
mem[1194] = 6'b101001;
mem[1195] = 6'b101010;
mem[1196] = 6'b000101;
mem[1197] = 6'b101010;
mem[1198] = 6'b111111;
mem[1199] = 6'b000101;
mem[1200] = 6'b000101;
mem[1201] = 6'b011010;
mem[1202] = 6'b000101;
mem[1203] = 6'b101010;
mem[1204] = 6'b111111;
mem[1205] = 6'b111111;
mem[1206] = 6'b111111;
mem[1207] = 6'b111111;
mem[1208] = 6'b111111;
mem[1209] = 6'b111111;
mem[1210] = 6'b111111;
mem[1211] = 6'b111111;
mem[1212] = 6'b111111;
mem[1213] = 6'b111111;
mem[1214] = 6'b111111;
mem[1215] = 6'b111111;
mem[1216] = 6'b111111;
mem[1217] = 6'b111111;
mem[1218] = 6'b111111;
mem[1219] = 6'b111111;
mem[1220] = 6'b111111;
mem[1221] = 6'b111111;
mem[1222] = 6'b111111;
mem[1223] = 6'b111111;
mem[1224] = 6'b111111;
mem[1225] = 6'b111111;
mem[1226] = 6'b111111;
mem[1227] = 6'b111111;
mem[1228] = 6'b101010;
mem[1229] = 6'b000101;
mem[1230] = 6'b000101;
mem[1231] = 6'b001001;
mem[1232] = 6'b011010;
mem[1233] = 6'b101010;
mem[1234] = 6'b101010;
mem[1235] = 6'b000101;
mem[1236] = 6'b111111;
mem[1237] = 6'b101010;
mem[1238] = 6'b000101;
mem[1239] = 6'b011010;
mem[1240] = 6'b000101;
mem[1241] = 6'b111010;
mem[1242] = 6'b101001;
mem[1243] = 6'b100100;
mem[1244] = 6'b000101;
mem[1245] = 6'b000101;
mem[1246] = 6'b101010;
mem[1247] = 6'b000101;
mem[1248] = 6'b000101;
mem[1249] = 6'b000101;
mem[1250] = 6'b101010;
mem[1251] = 6'b000101;
mem[1252] = 6'b101010;
mem[1253] = 6'b100101;
mem[1254] = 6'b100100;
mem[1255] = 6'b100100;
mem[1256] = 6'b101001;
mem[1257] = 6'b100100;
mem[1258] = 6'b101010;
mem[1259] = 6'b100100;
mem[1260] = 6'b100100;
mem[1261] = 6'b111111;
mem[1262] = 6'b000101;
mem[1263] = 6'b111111;
mem[1264] = 6'b101010;
mem[1265] = 6'b000101;
mem[1266] = 6'b000101;
mem[1267] = 6'b000101;
mem[1268] = 6'b111111;
mem[1269] = 6'b111111;
mem[1270] = 6'b111111;
mem[1271] = 6'b111111;
mem[1272] = 6'b111111;
mem[1273] = 6'b111111;
mem[1274] = 6'b111111;
mem[1275] = 6'b111111;
mem[1276] = 6'b111111;
mem[1277] = 6'b111111;
mem[1278] = 6'b111111;
mem[1279] = 6'b111111;
mem[1280] = 6'b111111;
mem[1281] = 6'b111111;
mem[1282] = 6'b111111;
mem[1283] = 6'b111111;
mem[1284] = 6'b111111;
mem[1285] = 6'b111111;
mem[1286] = 6'b111111;
mem[1287] = 6'b111111;
mem[1288] = 6'b111111;
mem[1289] = 6'b111111;
mem[1290] = 6'b111111;
mem[1291] = 6'b111111;
mem[1292] = 6'b011010;
mem[1293] = 6'b000101;
mem[1294] = 6'b000101;
mem[1295] = 6'b000101;
mem[1296] = 6'b000101;
mem[1297] = 6'b000101;
mem[1298] = 6'b101010;
mem[1299] = 6'b101010;
mem[1300] = 6'b001001;
mem[1301] = 6'b000101;
mem[1302] = 6'b011010;
mem[1303] = 6'b000101;
mem[1304] = 6'b101010;
mem[1305] = 6'b100100;
mem[1306] = 6'b100100;
mem[1307] = 6'b101010;
mem[1308] = 6'b000101;
mem[1309] = 6'b000101;
mem[1310] = 6'b101010;
mem[1311] = 6'b001001;
mem[1312] = 6'b000101;
mem[1313] = 6'b101010;
mem[1314] = 6'b111111;
mem[1315] = 6'b100100;
mem[1316] = 6'b100100;
mem[1317] = 6'b100100;
mem[1318] = 6'b111111;
mem[1319] = 6'b101010;
mem[1320] = 6'b101001;
mem[1321] = 6'b100100;
mem[1322] = 6'b100100;
mem[1323] = 6'b100100;
mem[1324] = 6'b100100;
mem[1325] = 6'b101010;
mem[1326] = 6'b111111;
mem[1327] = 6'b000101;
mem[1328] = 6'b000101;
mem[1329] = 6'b111111;
mem[1330] = 6'b001001;
mem[1331] = 6'b000101;
mem[1332] = 6'b101010;
mem[1333] = 6'b111111;
mem[1334] = 6'b111111;
mem[1335] = 6'b111111;
mem[1336] = 6'b111111;
mem[1337] = 6'b111111;
mem[1338] = 6'b111111;
mem[1339] = 6'b111111;
mem[1340] = 6'b111111;
mem[1341] = 6'b111111;
mem[1342] = 6'b111111;
mem[1343] = 6'b111111;
mem[1344] = 6'b111111;
mem[1345] = 6'b111111;
mem[1346] = 6'b111111;
mem[1347] = 6'b111111;
mem[1348] = 6'b111111;
mem[1349] = 6'b111111;
mem[1350] = 6'b111111;
mem[1351] = 6'b111111;
mem[1352] = 6'b111111;
mem[1353] = 6'b111111;
mem[1354] = 6'b111111;
mem[1355] = 6'b011001;
mem[1356] = 6'b101010;
mem[1357] = 6'b000101;
mem[1358] = 6'b000101;
mem[1359] = 6'b011010;
mem[1360] = 6'b000101;
mem[1361] = 6'b000101;
mem[1362] = 6'b101010;
mem[1363] = 6'b001001;
mem[1364] = 6'b011010;
mem[1365] = 6'b111111;
mem[1366] = 6'b000101;
mem[1367] = 6'b101010;
mem[1368] = 6'b100101;
mem[1369] = 6'b100100;
mem[1370] = 6'b100100;
mem[1371] = 6'b111111;
mem[1372] = 6'b011010;
mem[1373] = 6'b101010;
mem[1374] = 6'b011010;
mem[1375] = 6'b011010;
mem[1376] = 6'b000101;
mem[1377] = 6'b111111;
mem[1378] = 6'b100100;
mem[1379] = 6'b101001;
mem[1380] = 6'b100100;
mem[1381] = 6'b101010;
mem[1382] = 6'b000101;
mem[1383] = 6'b111111;
mem[1384] = 6'b000101;
mem[1385] = 6'b001001;
mem[1386] = 6'b111111;
mem[1387] = 6'b100100;
mem[1388] = 6'b101010;
mem[1389] = 6'b100100;
mem[1390] = 6'b100101;
mem[1391] = 6'b000101;
mem[1392] = 6'b000101;
mem[1393] = 6'b011010;
mem[1394] = 6'b000101;
mem[1395] = 6'b011010;
mem[1396] = 6'b011001;
mem[1397] = 6'b111111;
mem[1398] = 6'b111111;
mem[1399] = 6'b111111;
mem[1400] = 6'b111111;
mem[1401] = 6'b111111;
mem[1402] = 6'b111111;
mem[1403] = 6'b111111;
mem[1404] = 6'b111111;
mem[1405] = 6'b111111;
mem[1406] = 6'b111111;
mem[1407] = 6'b111111;
mem[1408] = 6'b111111;
mem[1409] = 6'b111111;
mem[1410] = 6'b111111;
mem[1411] = 6'b111111;
mem[1412] = 6'b111111;
mem[1413] = 6'b111111;
mem[1414] = 6'b111111;
mem[1415] = 6'b111111;
mem[1416] = 6'b111111;
mem[1417] = 6'b111111;
mem[1418] = 6'b111111;
mem[1419] = 6'b000101;
mem[1420] = 6'b000101;
mem[1421] = 6'b000101;
mem[1422] = 6'b011001;
mem[1423] = 6'b000101;
mem[1424] = 6'b111111;
mem[1425] = 6'b011010;
mem[1426] = 6'b001001;
mem[1427] = 6'b000101;
mem[1428] = 6'b000101;
mem[1429] = 6'b000101;
mem[1430] = 6'b111111;
mem[1431] = 6'b100100;
mem[1432] = 6'b101010;
mem[1433] = 6'b111111;
mem[1434] = 6'b100101;
mem[1435] = 6'b000101;
mem[1436] = 6'b101010;
mem[1437] = 6'b000101;
mem[1438] = 6'b101010;
mem[1439] = 6'b111111;
mem[1440] = 6'b001001;
mem[1441] = 6'b100100;
mem[1442] = 6'b100100;
mem[1443] = 6'b100100;
mem[1444] = 6'b111111;
mem[1445] = 6'b011010;
mem[1446] = 6'b011010;
mem[1447] = 6'b001001;
mem[1448] = 6'b000101;
mem[1449] = 6'b000101;
mem[1450] = 6'b011010;
mem[1451] = 6'b111111;
mem[1452] = 6'b100100;
mem[1453] = 6'b101001;
mem[1454] = 6'b101010;
mem[1455] = 6'b101010;
mem[1456] = 6'b111111;
mem[1457] = 6'b000101;
mem[1458] = 6'b000101;
mem[1459] = 6'b111111;
mem[1460] = 6'b000101;
mem[1461] = 6'b101010;
mem[1462] = 6'b111111;
mem[1463] = 6'b111111;
mem[1464] = 6'b111111;
mem[1465] = 6'b111111;
mem[1466] = 6'b111111;
mem[1467] = 6'b111111;
mem[1468] = 6'b111111;
mem[1469] = 6'b111111;
mem[1470] = 6'b111111;
mem[1471] = 6'b111111;
mem[1472] = 6'b111111;
mem[1473] = 6'b111111;
mem[1474] = 6'b111111;
mem[1475] = 6'b111111;
mem[1476] = 6'b111111;
mem[1477] = 6'b111111;
mem[1478] = 6'b111111;
mem[1479] = 6'b111111;
mem[1480] = 6'b111111;
mem[1481] = 6'b111111;
mem[1482] = 6'b011010;
mem[1483] = 6'b011010;
mem[1484] = 6'b111111;
mem[1485] = 6'b011010;
mem[1486] = 6'b000101;
mem[1487] = 6'b000101;
mem[1488] = 6'b000101;
mem[1489] = 6'b000101;
mem[1490] = 6'b111111;
mem[1491] = 6'b011010;
mem[1492] = 6'b000101;
mem[1493] = 6'b001001;
mem[1494] = 6'b100100;
mem[1495] = 6'b100100;
mem[1496] = 6'b100100;
mem[1497] = 6'b101001;
mem[1498] = 6'b100100;
mem[1499] = 6'b111111;
mem[1500] = 6'b011001;
mem[1501] = 6'b101010;
mem[1502] = 6'b000101;
mem[1503] = 6'b000101;
mem[1504] = 6'b101010;
mem[1505] = 6'b111111;
mem[1506] = 6'b100100;
mem[1507] = 6'b100100;
mem[1508] = 6'b000101;
mem[1509] = 6'b000101;
mem[1510] = 6'b001001;
mem[1511] = 6'b111111;
mem[1512] = 6'b000101;
mem[1513] = 6'b101010;
mem[1514] = 6'b000101;
mem[1515] = 6'b000101;
mem[1516] = 6'b100100;
mem[1517] = 6'b100100;
mem[1518] = 6'b101010;
mem[1519] = 6'b101010;
mem[1520] = 6'b001001;
mem[1521] = 6'b000101;
mem[1522] = 6'b000101;
mem[1523] = 6'b101010;
mem[1524] = 6'b101010;
mem[1525] = 6'b011010;
mem[1526] = 6'b111111;
mem[1527] = 6'b111111;
mem[1528] = 6'b111111;
mem[1529] = 6'b111111;
mem[1530] = 6'b111111;
mem[1531] = 6'b111111;
mem[1532] = 6'b111111;
mem[1533] = 6'b111111;
mem[1534] = 6'b111111;
mem[1535] = 6'b111111;
mem[1536] = 6'b111111;
mem[1537] = 6'b111111;
mem[1538] = 6'b111111;
mem[1539] = 6'b111111;
mem[1540] = 6'b111111;
mem[1541] = 6'b111111;
mem[1542] = 6'b111111;
mem[1543] = 6'b111111;
mem[1544] = 6'b111111;
mem[1545] = 6'b111111;
mem[1546] = 6'b000101;
mem[1547] = 6'b000101;
mem[1548] = 6'b000101;
mem[1549] = 6'b000101;
mem[1550] = 6'b001001;
mem[1551] = 6'b101010;
mem[1552] = 6'b000101;
mem[1553] = 6'b111111;
mem[1554] = 6'b000101;
mem[1555] = 6'b011010;
mem[1556] = 6'b111010;
mem[1557] = 6'b100100;
mem[1558] = 6'b111111;
mem[1559] = 6'b111111;
mem[1560] = 6'b100100;
mem[1561] = 6'b101001;
mem[1562] = 6'b101001;
mem[1563] = 6'b000101;
mem[1564] = 6'b000101;
mem[1565] = 6'b011010;
mem[1566] = 6'b000101;
mem[1567] = 6'b000101;
mem[1568] = 6'b101010;
mem[1569] = 6'b100100;
mem[1570] = 6'b101010;
mem[1571] = 6'b100100;
mem[1572] = 6'b000101;
mem[1573] = 6'b000101;
mem[1574] = 6'b101010;
mem[1575] = 6'b000101;
mem[1576] = 6'b000101;
mem[1577] = 6'b000101;
mem[1578] = 6'b101010;
mem[1579] = 6'b111111;
mem[1580] = 6'b100100;
mem[1581] = 6'b100100;
mem[1582] = 6'b100101;
mem[1583] = 6'b100100;
mem[1584] = 6'b000101;
mem[1585] = 6'b000101;
mem[1586] = 6'b101010;
mem[1587] = 6'b011010;
mem[1588] = 6'b000101;
mem[1589] = 6'b000101;
mem[1590] = 6'b111111;
mem[1591] = 6'b111111;
mem[1592] = 6'b111111;
mem[1593] = 6'b111111;
mem[1594] = 6'b111111;
mem[1595] = 6'b111111;
mem[1596] = 6'b111111;
mem[1597] = 6'b111111;
mem[1598] = 6'b111111;
mem[1599] = 6'b111111;
mem[1600] = 6'b111111;
mem[1601] = 6'b111111;
mem[1602] = 6'b111111;
mem[1603] = 6'b111111;
mem[1604] = 6'b111111;
mem[1605] = 6'b111111;
mem[1606] = 6'b111111;
mem[1607] = 6'b111111;
mem[1608] = 6'b111111;
mem[1609] = 6'b111111;
mem[1610] = 6'b000101;
mem[1611] = 6'b101010;
mem[1612] = 6'b000101;
mem[1613] = 6'b000101;
mem[1614] = 6'b101010;
mem[1615] = 6'b000101;
mem[1616] = 6'b101010;
mem[1617] = 6'b000101;
mem[1618] = 6'b000101;
mem[1619] = 6'b100100;
mem[1620] = 6'b101010;
mem[1621] = 6'b100100;
mem[1622] = 6'b001001;
mem[1623] = 6'b111111;
mem[1624] = 6'b100100;
mem[1625] = 6'b111111;
mem[1626] = 6'b100101;
mem[1627] = 6'b000101;
mem[1628] = 6'b000101;
mem[1629] = 6'b101111;
mem[1630] = 6'b111111;
mem[1631] = 6'b111111;
mem[1632] = 6'b100100;
mem[1633] = 6'b111111;
mem[1634] = 6'b101010;
mem[1635] = 6'b100100;
mem[1636] = 6'b100100;
mem[1637] = 6'b111010;
mem[1638] = 6'b001001;
mem[1639] = 6'b011010;
mem[1640] = 6'b111111;
mem[1641] = 6'b000101;
mem[1642] = 6'b001001;
mem[1643] = 6'b101010;
mem[1644] = 6'b101010;
mem[1645] = 6'b100100;
mem[1646] = 6'b100100;
mem[1647] = 6'b100100;
mem[1648] = 6'b000101;
mem[1649] = 6'b000101;
mem[1650] = 6'b101010;
mem[1651] = 6'b101110;
mem[1652] = 6'b000101;
mem[1653] = 6'b000101;
mem[1654] = 6'b011010;
mem[1655] = 6'b111111;
mem[1656] = 6'b111111;
mem[1657] = 6'b111111;
mem[1658] = 6'b111111;
mem[1659] = 6'b111111;
mem[1660] = 6'b111111;
mem[1661] = 6'b111111;
mem[1662] = 6'b111111;
mem[1663] = 6'b111111;
mem[1664] = 6'b111111;
mem[1665] = 6'b111111;
mem[1666] = 6'b111111;
mem[1667] = 6'b111111;
mem[1668] = 6'b111111;
mem[1669] = 6'b111111;
mem[1670] = 6'b111111;
mem[1671] = 6'b111111;
mem[1672] = 6'b111111;
mem[1673] = 6'b011010;
mem[1674] = 6'b000101;
mem[1675] = 6'b111111;
mem[1676] = 6'b001001;
mem[1677] = 6'b001001;
mem[1678] = 6'b101010;
mem[1679] = 6'b000101;
mem[1680] = 6'b000101;
mem[1681] = 6'b000101;
mem[1682] = 6'b000101;
mem[1683] = 6'b101010;
mem[1684] = 6'b100100;
mem[1685] = 6'b001001;
mem[1686] = 6'b000101;
mem[1687] = 6'b100100;
mem[1688] = 6'b111010;
mem[1689] = 6'b100100;
mem[1690] = 6'b101010;
mem[1691] = 6'b000101;
mem[1692] = 6'b101010;
mem[1693] = 6'b000101;
mem[1694] = 6'b000101;
mem[1695] = 6'b000101;
mem[1696] = 6'b100100;
mem[1697] = 6'b100101;
mem[1698] = 6'b101010;
mem[1699] = 6'b101010;
mem[1700] = 6'b100100;
mem[1701] = 6'b100101;
mem[1702] = 6'b000101;
mem[1703] = 6'b000101;
mem[1704] = 6'b000101;
mem[1705] = 6'b000101;
mem[1706] = 6'b000101;
mem[1707] = 6'b100100;
mem[1708] = 6'b100100;
mem[1709] = 6'b100100;
mem[1710] = 6'b100101;
mem[1711] = 6'b100100;
mem[1712] = 6'b111111;
mem[1713] = 6'b101010;
mem[1714] = 6'b011010;
mem[1715] = 6'b000101;
mem[1716] = 6'b101010;
mem[1717] = 6'b011010;
mem[1718] = 6'b000101;
mem[1719] = 6'b111111;
mem[1720] = 6'b111111;
mem[1721] = 6'b111111;
mem[1722] = 6'b111111;
mem[1723] = 6'b111111;
mem[1724] = 6'b111111;
mem[1725] = 6'b111111;
mem[1726] = 6'b111111;
mem[1727] = 6'b111111;
mem[1728] = 6'b111111;
mem[1729] = 6'b111111;
mem[1730] = 6'b111111;
mem[1731] = 6'b111111;
mem[1732] = 6'b111111;
mem[1733] = 6'b111111;
mem[1734] = 6'b111111;
mem[1735] = 6'b111111;
mem[1736] = 6'b111111;
mem[1737] = 6'b101111;
mem[1738] = 6'b001001;
mem[1739] = 6'b001001;
mem[1740] = 6'b000101;
mem[1741] = 6'b011010;
mem[1742] = 6'b011010;
mem[1743] = 6'b000101;
mem[1744] = 6'b011010;
mem[1745] = 6'b011010;
mem[1746] = 6'b111111;
mem[1747] = 6'b111010;
mem[1748] = 6'b011010;
mem[1749] = 6'b101010;
mem[1750] = 6'b101010;
mem[1751] = 6'b111111;
mem[1752] = 6'b100100;
mem[1753] = 6'b101001;
mem[1754] = 6'b101010;
mem[1755] = 6'b001001;
mem[1756] = 6'b011001;
mem[1757] = 6'b000101;
mem[1758] = 6'b101010;
mem[1759] = 6'b101010;
mem[1760] = 6'b100100;
mem[1761] = 6'b100100;
mem[1762] = 6'b100100;
mem[1763] = 6'b100100;
mem[1764] = 6'b101001;
mem[1765] = 6'b101010;
mem[1766] = 6'b000101;
mem[1767] = 6'b000101;
mem[1768] = 6'b111111;
mem[1769] = 6'b000101;
mem[1770] = 6'b101010;
mem[1771] = 6'b100100;
mem[1772] = 6'b100101;
mem[1773] = 6'b111111;
mem[1774] = 6'b100100;
mem[1775] = 6'b001001;
mem[1776] = 6'b000101;
mem[1777] = 6'b000101;
mem[1778] = 6'b101010;
mem[1779] = 6'b000101;
mem[1780] = 6'b001001;
mem[1781] = 6'b111111;
mem[1782] = 6'b011010;
mem[1783] = 6'b111111;
mem[1784] = 6'b111111;
mem[1785] = 6'b111111;
mem[1786] = 6'b111111;
mem[1787] = 6'b111111;
mem[1788] = 6'b111111;
mem[1789] = 6'b111111;
mem[1790] = 6'b111111;
mem[1791] = 6'b111111;
mem[1792] = 6'b111111;
mem[1793] = 6'b111111;
mem[1794] = 6'b111111;
mem[1795] = 6'b111111;
mem[1796] = 6'b111111;
mem[1797] = 6'b111111;
mem[1798] = 6'b111111;
mem[1799] = 6'b111111;
mem[1800] = 6'b111111;
mem[1801] = 6'b000101;
mem[1802] = 6'b000101;
mem[1803] = 6'b011010;
mem[1804] = 6'b111111;
mem[1805] = 6'b000101;
mem[1806] = 6'b011010;
mem[1807] = 6'b000101;
mem[1808] = 6'b000101;
mem[1809] = 6'b000101;
mem[1810] = 6'b000101;
mem[1811] = 6'b101010;
mem[1812] = 6'b000101;
mem[1813] = 6'b000101;
mem[1814] = 6'b111111;
mem[1815] = 6'b111010;
mem[1816] = 6'b100100;
mem[1817] = 6'b100100;
mem[1818] = 6'b011001;
mem[1819] = 6'b000101;
mem[1820] = 6'b001001;
mem[1821] = 6'b000101;
mem[1822] = 6'b000101;
mem[1823] = 6'b000101;
mem[1824] = 6'b001001;
mem[1825] = 6'b100100;
mem[1826] = 6'b100100;
mem[1827] = 6'b100100;
mem[1828] = 6'b111111;
mem[1829] = 6'b101010;
mem[1830] = 6'b001001;
mem[1831] = 6'b001001;
mem[1832] = 6'b000101;
mem[1833] = 6'b101010;
mem[1834] = 6'b101010;
mem[1835] = 6'b101010;
mem[1836] = 6'b101010;
mem[1837] = 6'b101010;
mem[1838] = 6'b101010;
mem[1839] = 6'b011010;
mem[1840] = 6'b111111;
mem[1841] = 6'b000101;
mem[1842] = 6'b101010;
mem[1843] = 6'b001001;
mem[1844] = 6'b001001;
mem[1845] = 6'b000101;
mem[1846] = 6'b000101;
mem[1847] = 6'b101010;
mem[1848] = 6'b111111;
mem[1849] = 6'b111111;
mem[1850] = 6'b111111;
mem[1851] = 6'b111111;
mem[1852] = 6'b111111;
mem[1853] = 6'b111111;
mem[1854] = 6'b111111;
mem[1855] = 6'b111111;
mem[1856] = 6'b111111;
mem[1857] = 6'b111111;
mem[1858] = 6'b111111;
mem[1859] = 6'b111111;
mem[1860] = 6'b111111;
mem[1861] = 6'b111111;
mem[1862] = 6'b111111;
mem[1863] = 6'b111111;
mem[1864] = 6'b111111;
mem[1865] = 6'b000101;
mem[1866] = 6'b000101;
mem[1867] = 6'b101010;
mem[1868] = 6'b000101;
mem[1869] = 6'b101010;
mem[1870] = 6'b111111;
mem[1871] = 6'b000101;
mem[1872] = 6'b011010;
mem[1873] = 6'b101010;
mem[1874] = 6'b011010;
mem[1875] = 6'b111111;
mem[1876] = 6'b000101;
mem[1877] = 6'b000101;
mem[1878] = 6'b100100;
mem[1879] = 6'b101001;
mem[1880] = 6'b100100;
mem[1881] = 6'b100100;
mem[1882] = 6'b011010;
mem[1883] = 6'b000101;
mem[1884] = 6'b000101;
mem[1885] = 6'b101010;
mem[1886] = 6'b000101;
mem[1887] = 6'b000101;
mem[1888] = 6'b000101;
mem[1889] = 6'b000101;
mem[1890] = 6'b011010;
mem[1891] = 6'b101010;
mem[1892] = 6'b011010;
mem[1893] = 6'b000101;
mem[1894] = 6'b111111;
mem[1895] = 6'b101010;
mem[1896] = 6'b001001;
mem[1897] = 6'b111111;
mem[1898] = 6'b100100;
mem[1899] = 6'b101010;
mem[1900] = 6'b100100;
mem[1901] = 6'b111111;
mem[1902] = 6'b000101;
mem[1903] = 6'b000101;
mem[1904] = 6'b001001;
mem[1905] = 6'b000101;
mem[1906] = 6'b101010;
mem[1907] = 6'b000101;
mem[1908] = 6'b000101;
mem[1909] = 6'b000101;
mem[1910] = 6'b000101;
mem[1911] = 6'b111111;
mem[1912] = 6'b111111;
mem[1913] = 6'b111111;
mem[1914] = 6'b111111;
mem[1915] = 6'b111111;
mem[1916] = 6'b111111;
mem[1917] = 6'b111111;
mem[1918] = 6'b111111;
mem[1919] = 6'b111111;
mem[1920] = 6'b111111;
mem[1921] = 6'b111111;
mem[1922] = 6'b111111;
mem[1923] = 6'b111111;
mem[1924] = 6'b111111;
mem[1925] = 6'b111111;
mem[1926] = 6'b111111;
mem[1927] = 6'b111111;
mem[1928] = 6'b111111;
mem[1929] = 6'b101010;
mem[1930] = 6'b000101;
mem[1931] = 6'b000101;
mem[1932] = 6'b000101;
mem[1933] = 6'b000101;
mem[1934] = 6'b000101;
mem[1935] = 6'b101010;
mem[1936] = 6'b000101;
mem[1937] = 6'b000101;
mem[1938] = 6'b000101;
mem[1939] = 6'b000101;
mem[1940] = 6'b000101;
mem[1941] = 6'b101010;
mem[1942] = 6'b101001;
mem[1943] = 6'b100100;
mem[1944] = 6'b100100;
mem[1945] = 6'b101010;
mem[1946] = 6'b111111;
mem[1947] = 6'b000101;
mem[1948] = 6'b000101;
mem[1949] = 6'b011010;
mem[1950] = 6'b011010;
mem[1951] = 6'b111111;
mem[1952] = 6'b111111;
mem[1953] = 6'b000101;
mem[1954] = 6'b001001;
mem[1955] = 6'b001001;
mem[1956] = 6'b000101;
mem[1957] = 6'b101010;
mem[1958] = 6'b000101;
mem[1959] = 6'b111111;
mem[1960] = 6'b100100;
mem[1961] = 6'b100100;
mem[1962] = 6'b101010;
mem[1963] = 6'b100100;
mem[1964] = 6'b101010;
mem[1965] = 6'b101010;
mem[1966] = 6'b000101;
mem[1967] = 6'b000101;
mem[1968] = 6'b101010;
mem[1969] = 6'b000101;
mem[1970] = 6'b011010;
mem[1971] = 6'b000101;
mem[1972] = 6'b000101;
mem[1973] = 6'b011010;
mem[1974] = 6'b000101;
mem[1975] = 6'b011010;
mem[1976] = 6'b111111;
mem[1977] = 6'b111111;
mem[1978] = 6'b111111;
mem[1979] = 6'b111111;
mem[1980] = 6'b111111;
mem[1981] = 6'b111111;
mem[1982] = 6'b111111;
mem[1983] = 6'b111111;
mem[1984] = 6'b111111;
mem[1985] = 6'b111111;
mem[1986] = 6'b111111;
mem[1987] = 6'b111111;
mem[1988] = 6'b111111;
mem[1989] = 6'b111111;
mem[1990] = 6'b111111;
mem[1991] = 6'b111111;
mem[1992] = 6'b000101;
mem[1993] = 6'b000101;
mem[1994] = 6'b011010;
mem[1995] = 6'b000101;
mem[1996] = 6'b000101;
mem[1997] = 6'b101010;
mem[1998] = 6'b101010;
mem[1999] = 6'b001001;
mem[2000] = 6'b000101;
mem[2001] = 6'b000101;
mem[2002] = 6'b101010;
mem[2003] = 6'b111111;
mem[2004] = 6'b000101;
mem[2005] = 6'b000101;
mem[2006] = 6'b101001;
mem[2007] = 6'b100100;
mem[2008] = 6'b101001;
mem[2009] = 6'b101010;
mem[2010] = 6'b000101;
mem[2011] = 6'b101010;
mem[2012] = 6'b000101;
mem[2013] = 6'b011010;
mem[2014] = 6'b000101;
mem[2015] = 6'b000101;
mem[2016] = 6'b000101;
mem[2017] = 6'b111111;
mem[2018] = 6'b101010;
mem[2019] = 6'b000101;
mem[2020] = 6'b000101;
mem[2021] = 6'b101010;
mem[2022] = 6'b111111;
mem[2023] = 6'b111111;
mem[2024] = 6'b100100;
mem[2025] = 6'b100100;
mem[2026] = 6'b111111;
mem[2027] = 6'b111111;
mem[2028] = 6'b000101;
mem[2029] = 6'b000101;
mem[2030] = 6'b000101;
mem[2031] = 6'b111111;
mem[2032] = 6'b001001;
mem[2033] = 6'b000101;
mem[2034] = 6'b111111;
mem[2035] = 6'b000101;
mem[2036] = 6'b011010;
mem[2037] = 6'b000101;
mem[2038] = 6'b000101;
mem[2039] = 6'b111111;
mem[2040] = 6'b111111;
mem[2041] = 6'b111111;
mem[2042] = 6'b111111;
mem[2043] = 6'b111111;
mem[2044] = 6'b111111;
mem[2045] = 6'b111111;
mem[2046] = 6'b111111;
mem[2047] = 6'b111111;
mem[2048] = 6'b111111;
mem[2049] = 6'b111111;
mem[2050] = 6'b111111;
mem[2051] = 6'b111111;
mem[2052] = 6'b111111;
mem[2053] = 6'b111111;
mem[2054] = 6'b111111;
mem[2055] = 6'b111111;
mem[2056] = 6'b111111;
mem[2057] = 6'b111111;
mem[2058] = 6'b001001;
mem[2059] = 6'b001001;
mem[2060] = 6'b001001;
mem[2061] = 6'b101010;
mem[2062] = 6'b000101;
mem[2063] = 6'b101010;
mem[2064] = 6'b101010;
mem[2065] = 6'b101010;
mem[2066] = 6'b000101;
mem[2067] = 6'b000101;
mem[2068] = 6'b000101;
mem[2069] = 6'b101010;
mem[2070] = 6'b100100;
mem[2071] = 6'b100101;
mem[2072] = 6'b100100;
mem[2073] = 6'b111111;
mem[2074] = 6'b011010;
mem[2075] = 6'b101010;
mem[2076] = 6'b000101;
mem[2077] = 6'b000101;
mem[2078] = 6'b101010;
mem[2079] = 6'b101010;
mem[2080] = 6'b111111;
mem[2081] = 6'b000101;
mem[2082] = 6'b000101;
mem[2083] = 6'b001001;
mem[2084] = 6'b000101;
mem[2085] = 6'b101010;
mem[2086] = 6'b101010;
mem[2087] = 6'b101010;
mem[2088] = 6'b101010;
mem[2089] = 6'b101010;
mem[2090] = 6'b000101;
mem[2091] = 6'b000101;
mem[2092] = 6'b011001;
mem[2093] = 6'b000101;
mem[2094] = 6'b101010;
mem[2095] = 6'b000101;
mem[2096] = 6'b011010;
mem[2097] = 6'b000101;
mem[2098] = 6'b101010;
mem[2099] = 6'b101010;
mem[2100] = 6'b000101;
mem[2101] = 6'b111111;
mem[2102] = 6'b111111;
mem[2103] = 6'b011010;
mem[2104] = 6'b111111;
mem[2105] = 6'b111111;
mem[2106] = 6'b111111;
mem[2107] = 6'b111111;
mem[2108] = 6'b111111;
mem[2109] = 6'b111111;
mem[2110] = 6'b111111;
mem[2111] = 6'b111111;
mem[2112] = 6'b111111;
mem[2113] = 6'b111111;
mem[2114] = 6'b111111;
mem[2115] = 6'b111111;
mem[2116] = 6'b111111;
mem[2117] = 6'b111111;
mem[2118] = 6'b111111;
mem[2119] = 6'b111111;
mem[2120] = 6'b101010;
mem[2121] = 6'b000101;
mem[2122] = 6'b101010;
mem[2123] = 6'b011001;
mem[2124] = 6'b000101;
mem[2125] = 6'b000101;
mem[2126] = 6'b000101;
mem[2127] = 6'b111111;
mem[2128] = 6'b101010;
mem[2129] = 6'b000101;
mem[2130] = 6'b111111;
mem[2131] = 6'b111111;
mem[2132] = 6'b001001;
mem[2133] = 6'b111111;
mem[2134] = 6'b101010;
mem[2135] = 6'b101001;
mem[2136] = 6'b111010;
mem[2137] = 6'b000101;
mem[2138] = 6'b000101;
mem[2139] = 6'b101111;
mem[2140] = 6'b000101;
mem[2141] = 6'b000101;
mem[2142] = 6'b101010;
mem[2143] = 6'b101010;
mem[2144] = 6'b101010;
mem[2145] = 6'b000101;
mem[2146] = 6'b000101;
mem[2147] = 6'b101010;
mem[2148] = 6'b111111;
mem[2149] = 6'b100100;
mem[2150] = 6'b100100;
mem[2151] = 6'b001001;
mem[2152] = 6'b000101;
mem[2153] = 6'b000101;
mem[2154] = 6'b000101;
mem[2155] = 6'b000101;
mem[2156] = 6'b011010;
mem[2157] = 6'b000101;
mem[2158] = 6'b101010;
mem[2159] = 6'b000101;
mem[2160] = 6'b000101;
mem[2161] = 6'b001001;
mem[2162] = 6'b000101;
mem[2163] = 6'b000101;
mem[2164] = 6'b111111;
mem[2165] = 6'b000101;
mem[2166] = 6'b000101;
mem[2167] = 6'b111111;
mem[2168] = 6'b111111;
mem[2169] = 6'b111111;
mem[2170] = 6'b111111;
mem[2171] = 6'b111111;
mem[2172] = 6'b111111;
mem[2173] = 6'b111111;
mem[2174] = 6'b111111;
mem[2175] = 6'b111111;
mem[2176] = 6'b111111;
mem[2177] = 6'b111111;
mem[2178] = 6'b111111;
mem[2179] = 6'b111111;
mem[2180] = 6'b111111;
mem[2181] = 6'b111111;
mem[2182] = 6'b111111;
mem[2183] = 6'b111111;
mem[2184] = 6'b111111;
mem[2185] = 6'b011010;
mem[2186] = 6'b111111;
mem[2187] = 6'b000101;
mem[2188] = 6'b000101;
mem[2189] = 6'b000101;
mem[2190] = 6'b000101;
mem[2191] = 6'b011010;
mem[2192] = 6'b000101;
mem[2193] = 6'b101010;
mem[2194] = 6'b001001;
mem[2195] = 6'b000101;
mem[2196] = 6'b000101;
mem[2197] = 6'b100100;
mem[2198] = 6'b111111;
mem[2199] = 6'b100100;
mem[2200] = 6'b111111;
mem[2201] = 6'b000101;
mem[2202] = 6'b000101;
mem[2203] = 6'b111111;
mem[2204] = 6'b000101;
mem[2205] = 6'b001001;
mem[2206] = 6'b000101;
mem[2207] = 6'b000101;
mem[2208] = 6'b111111;
mem[2209] = 6'b000101;
mem[2210] = 6'b001001;
mem[2211] = 6'b100100;
mem[2212] = 6'b100100;
mem[2213] = 6'b111111;
mem[2214] = 6'b101010;
mem[2215] = 6'b011010;
mem[2216] = 6'b001001;
mem[2217] = 6'b011010;
mem[2218] = 6'b101010;
mem[2219] = 6'b101010;
mem[2220] = 6'b000101;
mem[2221] = 6'b001001;
mem[2222] = 6'b101010;
mem[2223] = 6'b000101;
mem[2224] = 6'b000101;
mem[2225] = 6'b101110;
mem[2226] = 6'b000101;
mem[2227] = 6'b011010;
mem[2228] = 6'b011010;
mem[2229] = 6'b000101;
mem[2230] = 6'b000101;
mem[2231] = 6'b011010;
mem[2232] = 6'b111111;
mem[2233] = 6'b111111;
mem[2234] = 6'b111111;
mem[2235] = 6'b111111;
mem[2236] = 6'b111111;
mem[2237] = 6'b111111;
mem[2238] = 6'b111111;
mem[2239] = 6'b111111;
mem[2240] = 6'b111111;
mem[2241] = 6'b111111;
mem[2242] = 6'b111111;
mem[2243] = 6'b111111;
mem[2244] = 6'b111111;
mem[2245] = 6'b111111;
mem[2246] = 6'b111111;
mem[2247] = 6'b111111;
mem[2248] = 6'b111111;
mem[2249] = 6'b000101;
mem[2250] = 6'b000101;
mem[2251] = 6'b011010;
mem[2252] = 6'b101010;
mem[2253] = 6'b111111;
mem[2254] = 6'b001001;
mem[2255] = 6'b111111;
mem[2256] = 6'b000101;
mem[2257] = 6'b000101;
mem[2258] = 6'b011010;
mem[2259] = 6'b000101;
mem[2260] = 6'b000101;
mem[2261] = 6'b100100;
mem[2262] = 6'b100100;
mem[2263] = 6'b111111;
mem[2264] = 6'b000101;
mem[2265] = 6'b101010;
mem[2266] = 6'b101010;
mem[2267] = 6'b000101;
mem[2268] = 6'b000101;
mem[2269] = 6'b000101;
mem[2270] = 6'b111111;
mem[2271] = 6'b011010;
mem[2272] = 6'b000101;
mem[2273] = 6'b111111;
mem[2274] = 6'b100100;
mem[2275] = 6'b101010;
mem[2276] = 6'b111111;
mem[2277] = 6'b000101;
mem[2278] = 6'b000101;
mem[2279] = 6'b011010;
mem[2280] = 6'b000101;
mem[2281] = 6'b000101;
mem[2282] = 6'b000101;
mem[2283] = 6'b111111;
mem[2284] = 6'b001001;
mem[2285] = 6'b101010;
mem[2286] = 6'b001001;
mem[2287] = 6'b101010;
mem[2288] = 6'b101010;
mem[2289] = 6'b001001;
mem[2290] = 6'b000101;
mem[2291] = 6'b011010;
mem[2292] = 6'b101010;
mem[2293] = 6'b101010;
mem[2294] = 6'b001001;
mem[2295] = 6'b111111;
mem[2296] = 6'b111111;
mem[2297] = 6'b111111;
mem[2298] = 6'b111111;
mem[2299] = 6'b111111;
mem[2300] = 6'b111111;
mem[2301] = 6'b111111;
mem[2302] = 6'b111111;
mem[2303] = 6'b111111;
mem[2304] = 6'b111111;
mem[2305] = 6'b111111;
mem[2306] = 6'b111111;
mem[2307] = 6'b111111;
mem[2308] = 6'b111111;
mem[2309] = 6'b111111;
mem[2310] = 6'b111111;
mem[2311] = 6'b111111;
mem[2312] = 6'b111111;
mem[2313] = 6'b000101;
mem[2314] = 6'b000101;
mem[2315] = 6'b011010;
mem[2316] = 6'b000101;
mem[2317] = 6'b000101;
mem[2318] = 6'b000101;
mem[2319] = 6'b000101;
mem[2320] = 6'b011010;
mem[2321] = 6'b001001;
mem[2322] = 6'b001001;
mem[2323] = 6'b101010;
mem[2324] = 6'b111111;
mem[2325] = 6'b100100;
mem[2326] = 6'b100100;
mem[2327] = 6'b101010;
mem[2328] = 6'b101010;
mem[2329] = 6'b000101;
mem[2330] = 6'b111111;
mem[2331] = 6'b011010;
mem[2332] = 6'b101010;
mem[2333] = 6'b101010;
mem[2334] = 6'b000101;
mem[2335] = 6'b101010;
mem[2336] = 6'b100100;
mem[2337] = 6'b100100;
mem[2338] = 6'b101001;
mem[2339] = 6'b111111;
mem[2340] = 6'b001001;
mem[2341] = 6'b000101;
mem[2342] = 6'b000101;
mem[2343] = 6'b101010;
mem[2344] = 6'b001001;
mem[2345] = 6'b000101;
mem[2346] = 6'b101010;
mem[2347] = 6'b000101;
mem[2348] = 6'b000101;
mem[2349] = 6'b011010;
mem[2350] = 6'b000101;
mem[2351] = 6'b111111;
mem[2352] = 6'b000101;
mem[2353] = 6'b101010;
mem[2354] = 6'b011010;
mem[2355] = 6'b101010;
mem[2356] = 6'b101010;
mem[2357] = 6'b000101;
mem[2358] = 6'b000101;
mem[2359] = 6'b101010;
mem[2360] = 6'b111111;
mem[2361] = 6'b111111;
mem[2362] = 6'b111111;
mem[2363] = 6'b111111;
mem[2364] = 6'b111111;
mem[2365] = 6'b111111;
mem[2366] = 6'b111111;
mem[2367] = 6'b111111;
mem[2368] = 6'b111111;
mem[2369] = 6'b111111;
mem[2370] = 6'b111111;
mem[2371] = 6'b111111;
mem[2372] = 6'b111111;
mem[2373] = 6'b111111;
mem[2374] = 6'b111111;
mem[2375] = 6'b111111;
mem[2376] = 6'b111111;
mem[2377] = 6'b111111;
mem[2378] = 6'b101111;
mem[2379] = 6'b000101;
mem[2380] = 6'b000101;
mem[2381] = 6'b011010;
mem[2382] = 6'b000101;
mem[2383] = 6'b011010;
mem[2384] = 6'b000101;
mem[2385] = 6'b000101;
mem[2386] = 6'b111111;
mem[2387] = 6'b000101;
mem[2388] = 6'b000101;
mem[2389] = 6'b111010;
mem[2390] = 6'b100101;
mem[2391] = 6'b101010;
mem[2392] = 6'b101111;
mem[2393] = 6'b000101;
mem[2394] = 6'b101010;
mem[2395] = 6'b000101;
mem[2396] = 6'b000101;
mem[2397] = 6'b001001;
mem[2398] = 6'b000101;
mem[2399] = 6'b111111;
mem[2400] = 6'b100100;
mem[2401] = 6'b100100;
mem[2402] = 6'b111010;
mem[2403] = 6'b111010;
mem[2404] = 6'b100101;
mem[2405] = 6'b101010;
mem[2406] = 6'b100101;
mem[2407] = 6'b001001;
mem[2408] = 6'b000101;
mem[2409] = 6'b000101;
mem[2410] = 6'b101010;
mem[2411] = 6'b000101;
mem[2412] = 6'b000101;
mem[2413] = 6'b111111;
mem[2414] = 6'b111111;
mem[2415] = 6'b101010;
mem[2416] = 6'b101010;
mem[2417] = 6'b101010;
mem[2418] = 6'b000101;
mem[2419] = 6'b000101;
mem[2420] = 6'b111111;
mem[2421] = 6'b101010;
mem[2422] = 6'b000101;
mem[2423] = 6'b111111;
mem[2424] = 6'b111111;
mem[2425] = 6'b111111;
mem[2426] = 6'b111111;
mem[2427] = 6'b111111;
mem[2428] = 6'b111111;
mem[2429] = 6'b111111;
mem[2430] = 6'b111111;
mem[2431] = 6'b111111;
mem[2432] = 6'b111111;
mem[2433] = 6'b111111;
mem[2434] = 6'b111111;
mem[2435] = 6'b111111;
mem[2436] = 6'b111111;
mem[2437] = 6'b111111;
mem[2438] = 6'b111111;
mem[2439] = 6'b111111;
mem[2440] = 6'b111111;
mem[2441] = 6'b111111;
mem[2442] = 6'b000101;
mem[2443] = 6'b101010;
mem[2444] = 6'b001001;
mem[2445] = 6'b011001;
mem[2446] = 6'b011010;
mem[2447] = 6'b011010;
mem[2448] = 6'b001001;
mem[2449] = 6'b101010;
mem[2450] = 6'b000101;
mem[2451] = 6'b011010;
mem[2452] = 6'b100100;
mem[2453] = 6'b100100;
mem[2454] = 6'b111010;
mem[2455] = 6'b101001;
mem[2456] = 6'b000101;
mem[2457] = 6'b000101;
mem[2458] = 6'b111111;
mem[2459] = 6'b000101;
mem[2460] = 6'b000101;
mem[2461] = 6'b111111;
mem[2462] = 6'b100100;
mem[2463] = 6'b100100;
mem[2464] = 6'b100100;
mem[2465] = 6'b100100;
mem[2466] = 6'b101010;
mem[2467] = 6'b100100;
mem[2468] = 6'b100100;
mem[2469] = 6'b100100;
mem[2470] = 6'b100100;
mem[2471] = 6'b100100;
mem[2472] = 6'b100100;
mem[2473] = 6'b101010;
mem[2474] = 6'b001001;
mem[2475] = 6'b101010;
mem[2476] = 6'b111010;
mem[2477] = 6'b100100;
mem[2478] = 6'b000101;
mem[2479] = 6'b000101;
mem[2480] = 6'b001001;
mem[2481] = 6'b101010;
mem[2482] = 6'b000101;
mem[2483] = 6'b000101;
mem[2484] = 6'b101010;
mem[2485] = 6'b000101;
mem[2486] = 6'b101010;
mem[2487] = 6'b111111;
mem[2488] = 6'b111111;
mem[2489] = 6'b111111;
mem[2490] = 6'b111111;
mem[2491] = 6'b111111;
mem[2492] = 6'b111111;
mem[2493] = 6'b111111;
mem[2494] = 6'b111111;
mem[2495] = 6'b111111;
mem[2496] = 6'b111111;
mem[2497] = 6'b111111;
mem[2498] = 6'b111111;
mem[2499] = 6'b111111;
mem[2500] = 6'b111111;
mem[2501] = 6'b111111;
mem[2502] = 6'b111111;
mem[2503] = 6'b111111;
mem[2504] = 6'b111111;
mem[2505] = 6'b111111;
mem[2506] = 6'b000101;
mem[2507] = 6'b000101;
mem[2508] = 6'b101010;
mem[2509] = 6'b000101;
mem[2510] = 6'b101010;
mem[2511] = 6'b101010;
mem[2512] = 6'b011010;
mem[2513] = 6'b000101;
mem[2514] = 6'b000101;
mem[2515] = 6'b000101;
mem[2516] = 6'b101010;
mem[2517] = 6'b100100;
mem[2518] = 6'b101010;
mem[2519] = 6'b111111;
mem[2520] = 6'b000101;
mem[2521] = 6'b000101;
mem[2522] = 6'b101010;
mem[2523] = 6'b000101;
mem[2524] = 6'b000101;
mem[2525] = 6'b101010;
mem[2526] = 6'b100100;
mem[2527] = 6'b100100;
mem[2528] = 6'b100101;
mem[2529] = 6'b100100;
mem[2530] = 6'b100100;
mem[2531] = 6'b100100;
mem[2532] = 6'b100100;
mem[2533] = 6'b100101;
mem[2534] = 6'b100100;
mem[2535] = 6'b100100;
mem[2536] = 6'b101001;
mem[2537] = 6'b101010;
mem[2538] = 6'b101010;
mem[2539] = 6'b100100;
mem[2540] = 6'b100100;
mem[2541] = 6'b101010;
mem[2542] = 6'b000101;
mem[2543] = 6'b101010;
mem[2544] = 6'b000101;
mem[2545] = 6'b101010;
mem[2546] = 6'b101010;
mem[2547] = 6'b001001;
mem[2548] = 6'b000101;
mem[2549] = 6'b011010;
mem[2550] = 6'b111111;
mem[2551] = 6'b111111;
mem[2552] = 6'b111111;
mem[2553] = 6'b111111;
mem[2554] = 6'b111111;
mem[2555] = 6'b111111;
mem[2556] = 6'b111111;
mem[2557] = 6'b111111;
mem[2558] = 6'b111111;
mem[2559] = 6'b111111;
mem[2560] = 6'b111111;
mem[2561] = 6'b111111;
mem[2562] = 6'b111111;
mem[2563] = 6'b111111;
mem[2564] = 6'b111111;
mem[2565] = 6'b111111;
mem[2566] = 6'b111111;
mem[2567] = 6'b111111;
mem[2568] = 6'b111111;
mem[2569] = 6'b111111;
mem[2570] = 6'b101010;
mem[2571] = 6'b101010;
mem[2572] = 6'b000101;
mem[2573] = 6'b000101;
mem[2574] = 6'b000101;
mem[2575] = 6'b000101;
mem[2576] = 6'b000101;
mem[2577] = 6'b101010;
mem[2578] = 6'b001001;
mem[2579] = 6'b111111;
mem[2580] = 6'b101010;
mem[2581] = 6'b100100;
mem[2582] = 6'b100100;
mem[2583] = 6'b100100;
mem[2584] = 6'b011010;
mem[2585] = 6'b011001;
mem[2586] = 6'b101010;
mem[2587] = 6'b101010;
mem[2588] = 6'b101010;
mem[2589] = 6'b111010;
mem[2590] = 6'b100100;
mem[2591] = 6'b100101;
mem[2592] = 6'b101010;
mem[2593] = 6'b101010;
mem[2594] = 6'b101010;
mem[2595] = 6'b101010;
mem[2596] = 6'b111111;
mem[2597] = 6'b100100;
mem[2598] = 6'b101010;
mem[2599] = 6'b101010;
mem[2600] = 6'b100100;
mem[2601] = 6'b100100;
mem[2602] = 6'b101010;
mem[2603] = 6'b100100;
mem[2604] = 6'b100100;
mem[2605] = 6'b000101;
mem[2606] = 6'b000101;
mem[2607] = 6'b000101;
mem[2608] = 6'b101010;
mem[2609] = 6'b000101;
mem[2610] = 6'b000101;
mem[2611] = 6'b000101;
mem[2612] = 6'b000101;
mem[2613] = 6'b000101;
mem[2614] = 6'b111111;
mem[2615] = 6'b111111;
mem[2616] = 6'b111111;
mem[2617] = 6'b111111;
mem[2618] = 6'b111111;
mem[2619] = 6'b111111;
mem[2620] = 6'b111111;
mem[2621] = 6'b111111;
mem[2622] = 6'b111111;
mem[2623] = 6'b111111;
mem[2624] = 6'b111111;
mem[2625] = 6'b111111;
mem[2626] = 6'b111111;
mem[2627] = 6'b111111;
mem[2628] = 6'b111111;
mem[2629] = 6'b111111;
mem[2630] = 6'b111111;
mem[2631] = 6'b111111;
mem[2632] = 6'b111111;
mem[2633] = 6'b111111;
mem[2634] = 6'b111111;
mem[2635] = 6'b111111;
mem[2636] = 6'b000101;
mem[2637] = 6'b000101;
mem[2638] = 6'b101010;
mem[2639] = 6'b000101;
mem[2640] = 6'b000101;
mem[2641] = 6'b100100;
mem[2642] = 6'b100100;
mem[2643] = 6'b100100;
mem[2644] = 6'b100100;
mem[2645] = 6'b100100;
mem[2646] = 6'b100100;
mem[2647] = 6'b100100;
mem[2648] = 6'b100100;
mem[2649] = 6'b100100;
mem[2650] = 6'b000101;
mem[2651] = 6'b000101;
mem[2652] = 6'b100100;
mem[2653] = 6'b100100;
mem[2654] = 6'b000101;
mem[2655] = 6'b000101;
mem[2656] = 6'b000101;
mem[2657] = 6'b000101;
mem[2658] = 6'b000101;
mem[2659] = 6'b000101;
mem[2660] = 6'b111111;
mem[2661] = 6'b101010;
mem[2662] = 6'b100100;
mem[2663] = 6'b111111;
mem[2664] = 6'b100100;
mem[2665] = 6'b100100;
mem[2666] = 6'b100100;
mem[2667] = 6'b001001;
mem[2668] = 6'b101010;
mem[2669] = 6'b101111;
mem[2670] = 6'b000101;
mem[2671] = 6'b101010;
mem[2672] = 6'b001001;
mem[2673] = 6'b000101;
mem[2674] = 6'b111111;
mem[2675] = 6'b000101;
mem[2676] = 6'b001001;
mem[2677] = 6'b111111;
mem[2678] = 6'b111111;
mem[2679] = 6'b111111;
mem[2680] = 6'b111111;
mem[2681] = 6'b111111;
mem[2682] = 6'b111111;
mem[2683] = 6'b111111;
mem[2684] = 6'b111111;
mem[2685] = 6'b111111;
mem[2686] = 6'b111111;
mem[2687] = 6'b111111;
mem[2688] = 6'b111111;
mem[2689] = 6'b111111;
mem[2690] = 6'b111111;
mem[2691] = 6'b111111;
mem[2692] = 6'b111111;
mem[2693] = 6'b111111;
mem[2694] = 6'b111111;
mem[2695] = 6'b111111;
mem[2696] = 6'b111111;
mem[2697] = 6'b111111;
mem[2698] = 6'b111111;
mem[2699] = 6'b111111;
mem[2700] = 6'b000101;
mem[2701] = 6'b000101;
mem[2702] = 6'b000101;
mem[2703] = 6'b011010;
mem[2704] = 6'b101010;
mem[2705] = 6'b111111;
mem[2706] = 6'b111111;
mem[2707] = 6'b101010;
mem[2708] = 6'b011001;
mem[2709] = 6'b101010;
mem[2710] = 6'b111111;
mem[2711] = 6'b001001;
mem[2712] = 6'b111111;
mem[2713] = 6'b101010;
mem[2714] = 6'b000101;
mem[2715] = 6'b101010;
mem[2716] = 6'b111111;
mem[2717] = 6'b001001;
mem[2718] = 6'b101010;
mem[2719] = 6'b000101;
mem[2720] = 6'b000101;
mem[2721] = 6'b011010;
mem[2722] = 6'b011010;
mem[2723] = 6'b001001;
mem[2724] = 6'b111111;
mem[2725] = 6'b101110;
mem[2726] = 6'b000101;
mem[2727] = 6'b000101;
mem[2728] = 6'b001001;
mem[2729] = 6'b011010;
mem[2730] = 6'b001001;
mem[2731] = 6'b000101;
mem[2732] = 6'b001001;
mem[2733] = 6'b000101;
mem[2734] = 6'b000101;
mem[2735] = 6'b000101;
mem[2736] = 6'b000101;
mem[2737] = 6'b000101;
mem[2738] = 6'b101010;
mem[2739] = 6'b000101;
mem[2740] = 6'b000101;
mem[2741] = 6'b111111;
mem[2742] = 6'b111111;
mem[2743] = 6'b111111;
mem[2744] = 6'b111111;
mem[2745] = 6'b111111;
mem[2746] = 6'b111111;
mem[2747] = 6'b111111;
mem[2748] = 6'b111111;
mem[2749] = 6'b111111;
mem[2750] = 6'b111111;
mem[2751] = 6'b111111;
mem[2752] = 6'b111111;
mem[2753] = 6'b111111;
mem[2754] = 6'b111111;
mem[2755] = 6'b111111;
mem[2756] = 6'b111111;
mem[2757] = 6'b111111;
mem[2758] = 6'b111111;
mem[2759] = 6'b111111;
mem[2760] = 6'b111111;
mem[2761] = 6'b111111;
mem[2762] = 6'b111111;
mem[2763] = 6'b101010;
mem[2764] = 6'b000101;
mem[2765] = 6'b011010;
mem[2766] = 6'b000101;
mem[2767] = 6'b101010;
mem[2768] = 6'b011010;
mem[2769] = 6'b101010;
mem[2770] = 6'b000101;
mem[2771] = 6'b000101;
mem[2772] = 6'b111111;
mem[2773] = 6'b011001;
mem[2774] = 6'b000101;
mem[2775] = 6'b101010;
mem[2776] = 6'b111111;
mem[2777] = 6'b000101;
mem[2778] = 6'b000101;
mem[2779] = 6'b000101;
mem[2780] = 6'b000101;
mem[2781] = 6'b101010;
mem[2782] = 6'b000101;
mem[2783] = 6'b101010;
mem[2784] = 6'b011010;
mem[2785] = 6'b101010;
mem[2786] = 6'b011010;
mem[2787] = 6'b011010;
mem[2788] = 6'b000101;
mem[2789] = 6'b101010;
mem[2790] = 6'b000101;
mem[2791] = 6'b000101;
mem[2792] = 6'b101010;
mem[2793] = 6'b001001;
mem[2794] = 6'b000101;
mem[2795] = 6'b011001;
mem[2796] = 6'b000101;
mem[2797] = 6'b101010;
mem[2798] = 6'b000101;
mem[2799] = 6'b000101;
mem[2800] = 6'b000101;
mem[2801] = 6'b000101;
mem[2802] = 6'b111111;
mem[2803] = 6'b000101;
mem[2804] = 6'b000101;
mem[2805] = 6'b111111;
mem[2806] = 6'b111111;
mem[2807] = 6'b111111;
mem[2808] = 6'b111111;
mem[2809] = 6'b111111;
mem[2810] = 6'b111111;
mem[2811] = 6'b111111;
mem[2812] = 6'b111111;
mem[2813] = 6'b111111;
mem[2814] = 6'b111111;
mem[2815] = 6'b111111;
mem[2816] = 6'b111111;
mem[2817] = 6'b111111;
mem[2818] = 6'b111111;
mem[2819] = 6'b111111;
mem[2820] = 6'b111111;
mem[2821] = 6'b111111;
mem[2822] = 6'b111111;
mem[2823] = 6'b111111;
mem[2824] = 6'b111111;
mem[2825] = 6'b111111;
mem[2826] = 6'b111111;
mem[2827] = 6'b111111;
mem[2828] = 6'b001001;
mem[2829] = 6'b011010;
mem[2830] = 6'b000101;
mem[2831] = 6'b001001;
mem[2832] = 6'b111111;
mem[2833] = 6'b011010;
mem[2834] = 6'b000101;
mem[2835] = 6'b000101;
mem[2836] = 6'b101010;
mem[2837] = 6'b101010;
mem[2838] = 6'b101010;
mem[2839] = 6'b000101;
mem[2840] = 6'b000101;
mem[2841] = 6'b001001;
mem[2842] = 6'b000101;
mem[2843] = 6'b101010;
mem[2844] = 6'b011010;
mem[2845] = 6'b101010;
mem[2846] = 6'b001001;
mem[2847] = 6'b000101;
mem[2848] = 6'b000101;
mem[2849] = 6'b000101;
mem[2850] = 6'b000101;
mem[2851] = 6'b000101;
mem[2852] = 6'b111111;
mem[2853] = 6'b101010;
mem[2854] = 6'b000101;
mem[2855] = 6'b000101;
mem[2856] = 6'b101010;
mem[2857] = 6'b101010;
mem[2858] = 6'b001001;
mem[2859] = 6'b000101;
mem[2860] = 6'b000101;
mem[2861] = 6'b000101;
mem[2862] = 6'b011010;
mem[2863] = 6'b101010;
mem[2864] = 6'b101010;
mem[2865] = 6'b000101;
mem[2866] = 6'b000101;
mem[2867] = 6'b000101;
mem[2868] = 6'b111111;
mem[2869] = 6'b111111;
mem[2870] = 6'b111111;
mem[2871] = 6'b111111;
mem[2872] = 6'b111111;
mem[2873] = 6'b111111;
mem[2874] = 6'b111111;
mem[2875] = 6'b111111;
mem[2876] = 6'b111111;
mem[2877] = 6'b111111;
mem[2878] = 6'b111111;
mem[2879] = 6'b111111;
mem[2880] = 6'b111111;
mem[2881] = 6'b111111;
mem[2882] = 6'b111111;
mem[2883] = 6'b111111;
mem[2884] = 6'b111111;
mem[2885] = 6'b111111;
mem[2886] = 6'b111111;
mem[2887] = 6'b111111;
mem[2888] = 6'b111111;
mem[2889] = 6'b111111;
mem[2890] = 6'b111111;
mem[2891] = 6'b111111;
mem[2892] = 6'b111111;
mem[2893] = 6'b011010;
mem[2894] = 6'b000101;
mem[2895] = 6'b000101;
mem[2896] = 6'b000101;
mem[2897] = 6'b000101;
mem[2898] = 6'b101010;
mem[2899] = 6'b101010;
mem[2900] = 6'b000101;
mem[2901] = 6'b101010;
mem[2902] = 6'b000101;
mem[2903] = 6'b111111;
mem[2904] = 6'b011010;
mem[2905] = 6'b000101;
mem[2906] = 6'b111111;
mem[2907] = 6'b000101;
mem[2908] = 6'b011010;
mem[2909] = 6'b101010;
mem[2910] = 6'b001001;
mem[2911] = 6'b011010;
mem[2912] = 6'b000101;
mem[2913] = 6'b001001;
mem[2914] = 6'b101110;
mem[2915] = 6'b101010;
mem[2916] = 6'b000101;
mem[2917] = 6'b000101;
mem[2918] = 6'b101010;
mem[2919] = 6'b000101;
mem[2920] = 6'b000101;
mem[2921] = 6'b000101;
mem[2922] = 6'b101010;
mem[2923] = 6'b101010;
mem[2924] = 6'b000101;
mem[2925] = 6'b111111;
mem[2926] = 6'b001001;
mem[2927] = 6'b101010;
mem[2928] = 6'b001001;
mem[2929] = 6'b000101;
mem[2930] = 6'b011010;
mem[2931] = 6'b111111;
mem[2932] = 6'b111111;
mem[2933] = 6'b111111;
mem[2934] = 6'b111111;
mem[2935] = 6'b111111;
mem[2936] = 6'b111111;
mem[2937] = 6'b111111;
mem[2938] = 6'b111111;
mem[2939] = 6'b111111;
mem[2940] = 6'b111111;
mem[2941] = 6'b111111;
mem[2942] = 6'b111111;
mem[2943] = 6'b111111;
mem[2944] = 6'b111111;
mem[2945] = 6'b111111;
mem[2946] = 6'b111111;
mem[2947] = 6'b111111;
mem[2948] = 6'b111111;
mem[2949] = 6'b111111;
mem[2950] = 6'b111111;
mem[2951] = 6'b111111;
mem[2952] = 6'b111111;
mem[2953] = 6'b111111;
mem[2954] = 6'b111111;
mem[2955] = 6'b111111;
mem[2956] = 6'b111111;
mem[2957] = 6'b111111;
mem[2958] = 6'b000101;
mem[2959] = 6'b011010;
mem[2960] = 6'b111111;
mem[2961] = 6'b111111;
mem[2962] = 6'b011010;
mem[2963] = 6'b101010;
mem[2964] = 6'b000101;
mem[2965] = 6'b101010;
mem[2966] = 6'b011010;
mem[2967] = 6'b111111;
mem[2968] = 6'b000101;
mem[2969] = 6'b000101;
mem[2970] = 6'b001001;
mem[2971] = 6'b000101;
mem[2972] = 6'b111111;
mem[2973] = 6'b000101;
mem[2974] = 6'b000101;
mem[2975] = 6'b011010;
mem[2976] = 6'b000101;
mem[2977] = 6'b111111;
mem[2978] = 6'b000101;
mem[2979] = 6'b001001;
mem[2980] = 6'b000101;
mem[2981] = 6'b000101;
mem[2982] = 6'b111111;
mem[2983] = 6'b000101;
mem[2984] = 6'b000101;
mem[2985] = 6'b000101;
mem[2986] = 6'b101010;
mem[2987] = 6'b111111;
mem[2988] = 6'b000101;
mem[2989] = 6'b111111;
mem[2990] = 6'b000101;
mem[2991] = 6'b000101;
mem[2992] = 6'b001001;
mem[2993] = 6'b000101;
mem[2994] = 6'b111111;
mem[2995] = 6'b111111;
mem[2996] = 6'b111111;
mem[2997] = 6'b111111;
mem[2998] = 6'b111111;
mem[2999] = 6'b111111;
mem[3000] = 6'b111111;
mem[3001] = 6'b111111;
mem[3002] = 6'b111111;
mem[3003] = 6'b111111;
mem[3004] = 6'b111111;
mem[3005] = 6'b111111;
mem[3006] = 6'b111111;
mem[3007] = 6'b111111;
mem[3008] = 6'b111111;
mem[3009] = 6'b111111;
mem[3010] = 6'b111111;
mem[3011] = 6'b111111;
mem[3012] = 6'b111111;
mem[3013] = 6'b111111;
mem[3014] = 6'b111111;
mem[3015] = 6'b111111;
mem[3016] = 6'b111111;
mem[3017] = 6'b111111;
mem[3018] = 6'b111111;
mem[3019] = 6'b111111;
mem[3020] = 6'b111111;
mem[3021] = 6'b111111;
mem[3022] = 6'b111111;
mem[3023] = 6'b000101;
mem[3024] = 6'b101010;
mem[3025] = 6'b011010;
mem[3026] = 6'b000101;
mem[3027] = 6'b001001;
mem[3028] = 6'b000101;
mem[3029] = 6'b000101;
mem[3030] = 6'b000101;
mem[3031] = 6'b000101;
mem[3032] = 6'b011001;
mem[3033] = 6'b000101;
mem[3034] = 6'b101010;
mem[3035] = 6'b011010;
mem[3036] = 6'b000101;
mem[3037] = 6'b000101;
mem[3038] = 6'b000101;
mem[3039] = 6'b101110;
mem[3040] = 6'b000101;
mem[3041] = 6'b101010;
mem[3042] = 6'b000101;
mem[3043] = 6'b001001;
mem[3044] = 6'b001001;
mem[3045] = 6'b011001;
mem[3046] = 6'b101010;
mem[3047] = 6'b000101;
mem[3048] = 6'b000101;
mem[3049] = 6'b111111;
mem[3050] = 6'b000101;
mem[3051] = 6'b101010;
mem[3052] = 6'b000101;
mem[3053] = 6'b011010;
mem[3054] = 6'b000101;
mem[3055] = 6'b000101;
mem[3056] = 6'b001001;
mem[3057] = 6'b111111;
mem[3058] = 6'b111111;
mem[3059] = 6'b111111;
mem[3060] = 6'b111111;
mem[3061] = 6'b111111;
mem[3062] = 6'b111111;
mem[3063] = 6'b111111;
mem[3064] = 6'b111111;
mem[3065] = 6'b111111;
mem[3066] = 6'b111111;
mem[3067] = 6'b111111;
mem[3068] = 6'b111111;
mem[3069] = 6'b111111;
mem[3070] = 6'b111111;
mem[3071] = 6'b111111;
mem[3072] = 6'b111111;
mem[3073] = 6'b111111;
mem[3074] = 6'b111111;
mem[3075] = 6'b111111;
mem[3076] = 6'b111111;
mem[3077] = 6'b111111;
mem[3078] = 6'b111111;
mem[3079] = 6'b111111;
mem[3080] = 6'b111111;
mem[3081] = 6'b111111;
mem[3082] = 6'b111111;
mem[3083] = 6'b111111;
mem[3084] = 6'b111111;
mem[3085] = 6'b111111;
mem[3086] = 6'b111111;
mem[3087] = 6'b101010;
mem[3088] = 6'b011010;
mem[3089] = 6'b000101;
mem[3090] = 6'b001001;
mem[3091] = 6'b101010;
mem[3092] = 6'b001001;
mem[3093] = 6'b101010;
mem[3094] = 6'b000101;
mem[3095] = 6'b000101;
mem[3096] = 6'b000101;
mem[3097] = 6'b101010;
mem[3098] = 6'b000101;
mem[3099] = 6'b111111;
mem[3100] = 6'b101010;
mem[3101] = 6'b000101;
mem[3102] = 6'b011010;
mem[3103] = 6'b000101;
mem[3104] = 6'b011001;
mem[3105] = 6'b111111;
mem[3106] = 6'b000101;
mem[3107] = 6'b000101;
mem[3108] = 6'b011010;
mem[3109] = 6'b101010;
mem[3110] = 6'b101010;
mem[3111] = 6'b001001;
mem[3112] = 6'b011010;
mem[3113] = 6'b111111;
mem[3114] = 6'b001001;
mem[3115] = 6'b111111;
mem[3116] = 6'b000101;
mem[3117] = 6'b011010;
mem[3118] = 6'b101010;
mem[3119] = 6'b101010;
mem[3120] = 6'b111111;
mem[3121] = 6'b111111;
mem[3122] = 6'b111111;
mem[3123] = 6'b111111;
mem[3124] = 6'b111111;
mem[3125] = 6'b111111;
mem[3126] = 6'b111111;
mem[3127] = 6'b111111;
mem[3128] = 6'b111111;
mem[3129] = 6'b111111;
mem[3130] = 6'b111111;
mem[3131] = 6'b111111;
mem[3132] = 6'b111111;
mem[3133] = 6'b111111;
mem[3134] = 6'b111111;
mem[3135] = 6'b111111;
mem[3136] = 6'b111111;
mem[3137] = 6'b111111;
mem[3138] = 6'b111111;
mem[3139] = 6'b111111;
mem[3140] = 6'b111111;
mem[3141] = 6'b111111;
mem[3142] = 6'b111111;
mem[3143] = 6'b111111;
mem[3144] = 6'b111111;
mem[3145] = 6'b111111;
mem[3146] = 6'b111111;
mem[3147] = 6'b111111;
mem[3148] = 6'b111111;
mem[3149] = 6'b111111;
mem[3150] = 6'b111111;
mem[3151] = 6'b111111;
mem[3152] = 6'b101010;
mem[3153] = 6'b001001;
mem[3154] = 6'b011010;
mem[3155] = 6'b000101;
mem[3156] = 6'b000101;
mem[3157] = 6'b101010;
mem[3158] = 6'b101010;
mem[3159] = 6'b000101;
mem[3160] = 6'b111111;
mem[3161] = 6'b111111;
mem[3162] = 6'b000101;
mem[3163] = 6'b111111;
mem[3164] = 6'b011010;
mem[3165] = 6'b000101;
mem[3166] = 6'b111111;
mem[3167] = 6'b111111;
mem[3168] = 6'b000101;
mem[3169] = 6'b111111;
mem[3170] = 6'b000101;
mem[3171] = 6'b000101;
mem[3172] = 6'b101010;
mem[3173] = 6'b000101;
mem[3174] = 6'b000101;
mem[3175] = 6'b011010;
mem[3176] = 6'b000101;
mem[3177] = 6'b000101;
mem[3178] = 6'b000101;
mem[3179] = 6'b000101;
mem[3180] = 6'b101010;
mem[3181] = 6'b000101;
mem[3182] = 6'b101010;
mem[3183] = 6'b101010;
mem[3184] = 6'b111111;
mem[3185] = 6'b111111;
mem[3186] = 6'b111111;
mem[3187] = 6'b111111;
mem[3188] = 6'b111111;
mem[3189] = 6'b111111;
mem[3190] = 6'b111111;
mem[3191] = 6'b111111;
mem[3192] = 6'b111111;
mem[3193] = 6'b111111;
mem[3194] = 6'b111111;
mem[3195] = 6'b111111;
mem[3196] = 6'b111111;
mem[3197] = 6'b111111;
mem[3198] = 6'b111111;
mem[3199] = 6'b111111;
mem[3200] = 6'b111111;
mem[3201] = 6'b111111;
mem[3202] = 6'b111111;
mem[3203] = 6'b111111;
mem[3204] = 6'b111111;
mem[3205] = 6'b111111;
mem[3206] = 6'b111111;
mem[3207] = 6'b111111;
mem[3208] = 6'b111111;
mem[3209] = 6'b111111;
mem[3210] = 6'b111111;
mem[3211] = 6'b111111;
mem[3212] = 6'b111111;
mem[3213] = 6'b111111;
mem[3214] = 6'b111111;
mem[3215] = 6'b111111;
mem[3216] = 6'b111111;
mem[3217] = 6'b111111;
mem[3218] = 6'b001001;
mem[3219] = 6'b000101;
mem[3220] = 6'b000101;
mem[3221] = 6'b000101;
mem[3222] = 6'b000101;
mem[3223] = 6'b011010;
mem[3224] = 6'b000101;
mem[3225] = 6'b000101;
mem[3226] = 6'b000101;
mem[3227] = 6'b000101;
mem[3228] = 6'b001001;
mem[3229] = 6'b000101;
mem[3230] = 6'b000101;
mem[3231] = 6'b000101;
mem[3232] = 6'b101010;
mem[3233] = 6'b101010;
mem[3234] = 6'b000101;
mem[3235] = 6'b001001;
mem[3236] = 6'b111111;
mem[3237] = 6'b000101;
mem[3238] = 6'b000101;
mem[3239] = 6'b011010;
mem[3240] = 6'b101010;
mem[3241] = 6'b001001;
mem[3242] = 6'b000101;
mem[3243] = 6'b000101;
mem[3244] = 6'b101010;
mem[3245] = 6'b000101;
mem[3246] = 6'b111111;
mem[3247] = 6'b111111;
mem[3248] = 6'b111111;
mem[3249] = 6'b111111;
mem[3250] = 6'b111111;
mem[3251] = 6'b111111;
mem[3252] = 6'b111111;
mem[3253] = 6'b111111;
mem[3254] = 6'b111111;
mem[3255] = 6'b111111;
mem[3256] = 6'b111111;
mem[3257] = 6'b111111;
mem[3258] = 6'b111111;
mem[3259] = 6'b111111;
mem[3260] = 6'b111111;
mem[3261] = 6'b111111;
mem[3262] = 6'b111111;
mem[3263] = 6'b111111;
mem[3264] = 6'b111111;
mem[3265] = 6'b111111;
mem[3266] = 6'b111111;
mem[3267] = 6'b111111;
mem[3268] = 6'b111111;
mem[3269] = 6'b111111;
mem[3270] = 6'b111111;
mem[3271] = 6'b111111;
mem[3272] = 6'b111111;
mem[3273] = 6'b111111;
mem[3274] = 6'b111111;
mem[3275] = 6'b111111;
mem[3276] = 6'b111111;
mem[3277] = 6'b111111;
mem[3278] = 6'b111111;
mem[3279] = 6'b111111;
mem[3280] = 6'b111111;
mem[3281] = 6'b111111;
mem[3282] = 6'b111111;
mem[3283] = 6'b101010;
mem[3284] = 6'b101010;
mem[3285] = 6'b000101;
mem[3286] = 6'b011010;
mem[3287] = 6'b011010;
mem[3288] = 6'b101010;
mem[3289] = 6'b011010;
mem[3290] = 6'b000101;
mem[3291] = 6'b000101;
mem[3292] = 6'b000101;
mem[3293] = 6'b111111;
mem[3294] = 6'b111111;
mem[3295] = 6'b000101;
mem[3296] = 6'b111111;
mem[3297] = 6'b101010;
mem[3298] = 6'b000101;
mem[3299] = 6'b000101;
mem[3300] = 6'b101010;
mem[3301] = 6'b101010;
mem[3302] = 6'b001001;
mem[3303] = 6'b001001;
mem[3304] = 6'b011010;
mem[3305] = 6'b000101;
mem[3306] = 6'b101010;
mem[3307] = 6'b101010;
mem[3308] = 6'b011010;
mem[3309] = 6'b111111;
mem[3310] = 6'b111111;
mem[3311] = 6'b111111;
mem[3312] = 6'b111111;
mem[3313] = 6'b111111;
mem[3314] = 6'b111111;
mem[3315] = 6'b111111;
mem[3316] = 6'b111111;
mem[3317] = 6'b111111;
mem[3318] = 6'b111111;
mem[3319] = 6'b111111;
mem[3320] = 6'b111111;
mem[3321] = 6'b111111;
mem[3322] = 6'b111111;
mem[3323] = 6'b111111;
mem[3324] = 6'b111111;
mem[3325] = 6'b111111;
mem[3326] = 6'b111111;
mem[3327] = 6'b111111;
mem[3328] = 6'b111111;
mem[3329] = 6'b111111;
mem[3330] = 6'b111111;
mem[3331] = 6'b111111;
mem[3332] = 6'b111111;
mem[3333] = 6'b111111;
mem[3334] = 6'b111111;
mem[3335] = 6'b111111;
mem[3336] = 6'b111111;
mem[3337] = 6'b111111;
mem[3338] = 6'b111111;
mem[3339] = 6'b111111;
mem[3340] = 6'b111111;
mem[3341] = 6'b111111;
mem[3342] = 6'b111111;
mem[3343] = 6'b111111;
mem[3344] = 6'b111111;
mem[3345] = 6'b111111;
mem[3346] = 6'b111111;
mem[3347] = 6'b111111;
mem[3348] = 6'b111111;
mem[3349] = 6'b111111;
mem[3350] = 6'b000101;
mem[3351] = 6'b000101;
mem[3352] = 6'b000101;
mem[3353] = 6'b000101;
mem[3354] = 6'b101010;
mem[3355] = 6'b101010;
mem[3356] = 6'b101010;
mem[3357] = 6'b000101;
mem[3358] = 6'b011010;
mem[3359] = 6'b011010;
mem[3360] = 6'b111111;
mem[3361] = 6'b000101;
mem[3362] = 6'b111111;
mem[3363] = 6'b101010;
mem[3364] = 6'b111111;
mem[3365] = 6'b101010;
mem[3366] = 6'b011010;
mem[3367] = 6'b000101;
mem[3368] = 6'b101010;
mem[3369] = 6'b000101;
mem[3370] = 6'b000101;
mem[3371] = 6'b111111;
mem[3372] = 6'b111111;
mem[3373] = 6'b111111;
mem[3374] = 6'b111111;
mem[3375] = 6'b111111;
mem[3376] = 6'b111111;
mem[3377] = 6'b111111;
mem[3378] = 6'b111111;
mem[3379] = 6'b111111;
mem[3380] = 6'b111111;
mem[3381] = 6'b111111;
mem[3382] = 6'b111111;
mem[3383] = 6'b111111;
mem[3384] = 6'b111111;
mem[3385] = 6'b111111;
mem[3386] = 6'b111111;
mem[3387] = 6'b111111;
mem[3388] = 6'b111111;
mem[3389] = 6'b111111;
mem[3390] = 6'b111111;
mem[3391] = 6'b111111;
mem[3392] = 6'b111111;
mem[3393] = 6'b111111;
mem[3394] = 6'b111111;
mem[3395] = 6'b111111;
mem[3396] = 6'b111111;
mem[3397] = 6'b111111;
mem[3398] = 6'b111111;
mem[3399] = 6'b111111;
mem[3400] = 6'b111111;
mem[3401] = 6'b111111;
mem[3402] = 6'b111111;
mem[3403] = 6'b111111;
mem[3404] = 6'b111111;
mem[3405] = 6'b111111;
mem[3406] = 6'b111111;
mem[3407] = 6'b111111;
mem[3408] = 6'b111111;
mem[3409] = 6'b111111;
mem[3410] = 6'b111111;
mem[3411] = 6'b111111;
mem[3412] = 6'b111111;
mem[3413] = 6'b111111;
mem[3414] = 6'b111111;
mem[3415] = 6'b111111;
mem[3416] = 6'b000101;
mem[3417] = 6'b000101;
mem[3418] = 6'b101010;
mem[3419] = 6'b000101;
mem[3420] = 6'b111111;
mem[3421] = 6'b011010;
mem[3422] = 6'b101010;
mem[3423] = 6'b000101;
mem[3424] = 6'b000101;
mem[3425] = 6'b111111;
mem[3426] = 6'b000101;
mem[3427] = 6'b000101;
mem[3428] = 6'b111111;
mem[3429] = 6'b000101;
mem[3430] = 6'b101010;
mem[3431] = 6'b000101;
mem[3432] = 6'b011010;
mem[3433] = 6'b111111;
mem[3434] = 6'b111111;
mem[3435] = 6'b111111;
mem[3436] = 6'b111111;
mem[3437] = 6'b111111;
mem[3438] = 6'b111111;
mem[3439] = 6'b111111;
mem[3440] = 6'b111111;
mem[3441] = 6'b111111;
mem[3442] = 6'b111111;
mem[3443] = 6'b111111;
mem[3444] = 6'b111111;
mem[3445] = 6'b111111;
mem[3446] = 6'b111111;
mem[3447] = 6'b111111;
mem[3448] = 6'b111111;
mem[3449] = 6'b111111;
mem[3450] = 6'b111111;
mem[3451] = 6'b111111;
mem[3452] = 6'b111111;
mem[3453] = 6'b111111;
mem[3454] = 6'b111111;
mem[3455] = 6'b111111;
mem[3456] = 6'b111111;
mem[3457] = 6'b111111;
mem[3458] = 6'b111111;
mem[3459] = 6'b111111;
mem[3460] = 6'b111111;
mem[3461] = 6'b111111;
mem[3462] = 6'b111111;
mem[3463] = 6'b111111;
mem[3464] = 6'b111111;
mem[3465] = 6'b111111;
mem[3466] = 6'b111111;
mem[3467] = 6'b111111;
mem[3468] = 6'b111111;
mem[3469] = 6'b111111;
mem[3470] = 6'b111111;
mem[3471] = 6'b111111;
mem[3472] = 6'b111111;
mem[3473] = 6'b111111;
mem[3474] = 6'b111111;
mem[3475] = 6'b111111;
mem[3476] = 6'b111111;
mem[3477] = 6'b111111;
mem[3478] = 6'b111111;
mem[3479] = 6'b111111;
mem[3480] = 6'b111111;
mem[3481] = 6'b111111;
mem[3482] = 6'b011010;
mem[3483] = 6'b101010;
mem[3484] = 6'b011010;
mem[3485] = 6'b000101;
mem[3486] = 6'b101010;
mem[3487] = 6'b000101;
mem[3488] = 6'b000101;
mem[3489] = 6'b111111;
mem[3490] = 6'b000101;
mem[3491] = 6'b000101;
mem[3492] = 6'b111111;
mem[3493] = 6'b000101;
mem[3494] = 6'b111111;
mem[3495] = 6'b111111;
mem[3496] = 6'b111111;
mem[3497] = 6'b111111;
mem[3498] = 6'b111111;
mem[3499] = 6'b111111;
mem[3500] = 6'b111111;
mem[3501] = 6'b111111;
mem[3502] = 6'b111111;
mem[3503] = 6'b111111;
mem[3504] = 6'b111111;
mem[3505] = 6'b111111;
mem[3506] = 6'b111111;
mem[3507] = 6'b111111;
mem[3508] = 6'b111111;
mem[3509] = 6'b111111;
mem[3510] = 6'b111111;
mem[3511] = 6'b111111;
mem[3512] = 6'b111111;
mem[3513] = 6'b111111;
mem[3514] = 6'b111111;
mem[3515] = 6'b111111;
mem[3516] = 6'b111111;
mem[3517] = 6'b111111;
mem[3518] = 6'b111111;
mem[3519] = 6'b111111;
mem[3520] = 6'b111111;
mem[3521] = 6'b111111;
mem[3522] = 6'b111111;
mem[3523] = 6'b111111;
mem[3524] = 6'b111111;
mem[3525] = 6'b111111;
mem[3526] = 6'b111111;
mem[3527] = 6'b111111;
mem[3528] = 6'b111111;
mem[3529] = 6'b111111;
mem[3530] = 6'b111111;
mem[3531] = 6'b111111;
mem[3532] = 6'b111111;
mem[3533] = 6'b111111;
mem[3534] = 6'b111111;
mem[3535] = 6'b111111;
mem[3536] = 6'b111111;
mem[3537] = 6'b111111;
mem[3538] = 6'b111111;
mem[3539] = 6'b111111;
mem[3540] = 6'b111111;
mem[3541] = 6'b111111;
mem[3542] = 6'b111111;
mem[3543] = 6'b111111;
mem[3544] = 6'b111111;
mem[3545] = 6'b111111;
mem[3546] = 6'b111111;
mem[3547] = 6'b111111;
mem[3548] = 6'b111111;
mem[3549] = 6'b111111;
mem[3550] = 6'b111111;
mem[3551] = 6'b101010;
mem[3552] = 6'b111111;
mem[3553] = 6'b011010;
mem[3554] = 6'b111111;
mem[3555] = 6'b111111;
mem[3556] = 6'b111111;
mem[3557] = 6'b111111;
mem[3558] = 6'b111111;
mem[3559] = 6'b111111;
mem[3560] = 6'b111111;
mem[3561] = 6'b111111;
mem[3562] = 6'b111111;
mem[3563] = 6'b111111;
mem[3564] = 6'b111111;
mem[3565] = 6'b111111;
mem[3566] = 6'b111111;
mem[3567] = 6'b111111;
mem[3568] = 6'b111111;
mem[3569] = 6'b111111;
mem[3570] = 6'b111111;
mem[3571] = 6'b111111;
mem[3572] = 6'b111111;
mem[3573] = 6'b111111;
mem[3574] = 6'b111111;
mem[3575] = 6'b111111;
mem[3576] = 6'b111111;
mem[3577] = 6'b111111;
mem[3578] = 6'b111111;
mem[3579] = 6'b111111;
mem[3580] = 6'b111111;
mem[3581] = 6'b111111;
mem[3582] = 6'b111111;
mem[3583] = 6'b111111;
mem[3584] = 6'b111111;
mem[3585] = 6'b111111;
mem[3586] = 6'b111111;
mem[3587] = 6'b111111;
mem[3588] = 6'b111111;
mem[3589] = 6'b111111;
mem[3590] = 6'b111111;
mem[3591] = 6'b111111;
mem[3592] = 6'b111111;
mem[3593] = 6'b111111;
mem[3594] = 6'b111111;
mem[3595] = 6'b111111;
mem[3596] = 6'b111111;
mem[3597] = 6'b111111;
mem[3598] = 6'b111111;
mem[3599] = 6'b111111;
mem[3600] = 6'b111111;
mem[3601] = 6'b111111;
mem[3602] = 6'b111111;
mem[3603] = 6'b111111;
mem[3604] = 6'b111111;
mem[3605] = 6'b111111;
mem[3606] = 6'b111111;
mem[3607] = 6'b111111;
mem[3608] = 6'b111111;
mem[3609] = 6'b111111;
mem[3610] = 6'b111111;
mem[3611] = 6'b111111;
mem[3612] = 6'b111111;
mem[3613] = 6'b111111;
mem[3614] = 6'b111111;
mem[3615] = 6'b111111;
mem[3616] = 6'b111111;
mem[3617] = 6'b111111;
mem[3618] = 6'b111111;
mem[3619] = 6'b111111;
mem[3620] = 6'b111111;
mem[3621] = 6'b111111;
mem[3622] = 6'b111111;
mem[3623] = 6'b111111;
mem[3624] = 6'b111111;
mem[3625] = 6'b111111;
mem[3626] = 6'b111111;
mem[3627] = 6'b111111;
mem[3628] = 6'b111111;
mem[3629] = 6'b111111;
mem[3630] = 6'b111111;
mem[3631] = 6'b111111;
mem[3632] = 6'b111111;
mem[3633] = 6'b111111;
mem[3634] = 6'b111111;
mem[3635] = 6'b111111;
mem[3636] = 6'b111111;
mem[3637] = 6'b111111;
mem[3638] = 6'b111111;
mem[3639] = 6'b111111;
mem[3640] = 6'b111111;
mem[3641] = 6'b111111;
mem[3642] = 6'b111111;
mem[3643] = 6'b111111;
mem[3644] = 6'b111111;
mem[3645] = 6'b111111;
mem[3646] = 6'b111111;
mem[3647] = 6'b111111;
mem[3648] = 6'b111111;
mem[3649] = 6'b111111;
mem[3650] = 6'b111111;
mem[3651] = 6'b111111;
mem[3652] = 6'b111111;
mem[3653] = 6'b111111;
mem[3654] = 6'b111111;
mem[3655] = 6'b111111;
mem[3656] = 6'b111111;
mem[3657] = 6'b111111;
mem[3658] = 6'b111111;
mem[3659] = 6'b111111;
mem[3660] = 6'b111111;
mem[3661] = 6'b111111;
mem[3662] = 6'b111111;
mem[3663] = 6'b111111;
mem[3664] = 6'b111111;
mem[3665] = 6'b111111;
mem[3666] = 6'b111111;
mem[3667] = 6'b111111;
mem[3668] = 6'b111111;
mem[3669] = 6'b111111;
mem[3670] = 6'b111111;
mem[3671] = 6'b111111;
mem[3672] = 6'b111111;
mem[3673] = 6'b111111;
mem[3674] = 6'b111111;
mem[3675] = 6'b111111;
mem[3676] = 6'b111111;
mem[3677] = 6'b111111;
mem[3678] = 6'b111111;
mem[3679] = 6'b111111;
mem[3680] = 6'b111111;
mem[3681] = 6'b111111;
mem[3682] = 6'b111111;
mem[3683] = 6'b111111;
mem[3684] = 6'b111111;
mem[3685] = 6'b111111;
mem[3686] = 6'b111111;
mem[3687] = 6'b111111;
mem[3688] = 6'b111111;
mem[3689] = 6'b111111;
mem[3690] = 6'b111111;
mem[3691] = 6'b111111;
mem[3692] = 6'b111111;
mem[3693] = 6'b111111;
mem[3694] = 6'b111111;
mem[3695] = 6'b111111;
mem[3696] = 6'b111111;
mem[3697] = 6'b111111;
mem[3698] = 6'b111111;
mem[3699] = 6'b111111;
mem[3700] = 6'b111111;
mem[3701] = 6'b111111;
mem[3702] = 6'b111111;
mem[3703] = 6'b111111;
mem[3704] = 6'b111111;
mem[3705] = 6'b111111;
mem[3706] = 6'b111111;
mem[3707] = 6'b111111;
mem[3708] = 6'b111111;
mem[3709] = 6'b111111;
mem[3710] = 6'b111111;
mem[3711] = 6'b111111;
mem[3712] = 6'b111111;
mem[3713] = 6'b111111;
mem[3714] = 6'b111111;
mem[3715] = 6'b111111;
mem[3716] = 6'b111111;
mem[3717] = 6'b111111;
mem[3718] = 6'b111111;
mem[3719] = 6'b111111;
mem[3720] = 6'b111111;
mem[3721] = 6'b111111;
mem[3722] = 6'b111111;
mem[3723] = 6'b111111;
mem[3724] = 6'b111111;
mem[3725] = 6'b111111;
mem[3726] = 6'b111111;
mem[3727] = 6'b111111;
mem[3728] = 6'b111111;
mem[3729] = 6'b111111;
mem[3730] = 6'b111111;
mem[3731] = 6'b111111;
mem[3732] = 6'b111111;
mem[3733] = 6'b111111;
mem[3734] = 6'b111111;
mem[3735] = 6'b111111;
mem[3736] = 6'b111111;
mem[3737] = 6'b111111;
mem[3738] = 6'b111111;
mem[3739] = 6'b111111;
mem[3740] = 6'b111111;
mem[3741] = 6'b111111;
mem[3742] = 6'b111111;
mem[3743] = 6'b111111;
mem[3744] = 6'b111111;
mem[3745] = 6'b111111;
mem[3746] = 6'b111111;
mem[3747] = 6'b111111;
mem[3748] = 6'b111111;
mem[3749] = 6'b111111;
mem[3750] = 6'b111111;
mem[3751] = 6'b111111;
mem[3752] = 6'b111111;
mem[3753] = 6'b111111;
mem[3754] = 6'b111111;
mem[3755] = 6'b111111;
mem[3756] = 6'b111111;
mem[3757] = 6'b111111;
mem[3758] = 6'b111111;
mem[3759] = 6'b111111;
mem[3760] = 6'b111111;
mem[3761] = 6'b111111;
mem[3762] = 6'b111111;
mem[3763] = 6'b111111;
mem[3764] = 6'b111111;
mem[3765] = 6'b111111;
mem[3766] = 6'b111111;
mem[3767] = 6'b111111;
mem[3768] = 6'b111111;
mem[3769] = 6'b111111;
mem[3770] = 6'b111111;
mem[3771] = 6'b111111;
mem[3772] = 6'b111111;
mem[3773] = 6'b111111;
mem[3774] = 6'b111111;
mem[3775] = 6'b111111;
mem[3776] = 6'b111111;
mem[3777] = 6'b111111;
mem[3778] = 6'b111111;
mem[3779] = 6'b111111;
mem[3780] = 6'b111111;
mem[3781] = 6'b111111;
mem[3782] = 6'b111111;
mem[3783] = 6'b111111;
mem[3784] = 6'b111111;
mem[3785] = 6'b111111;
mem[3786] = 6'b111111;
mem[3787] = 6'b111111;
mem[3788] = 6'b111111;
mem[3789] = 6'b111111;
mem[3790] = 6'b111111;
mem[3791] = 6'b111111;
mem[3792] = 6'b111111;
mem[3793] = 6'b111111;
mem[3794] = 6'b111111;
mem[3795] = 6'b111111;
mem[3796] = 6'b111111;
mem[3797] = 6'b111111;
mem[3798] = 6'b111111;
mem[3799] = 6'b111111;
mem[3800] = 6'b111111;
mem[3801] = 6'b111111;
mem[3802] = 6'b111111;
mem[3803] = 6'b111111;
mem[3804] = 6'b111111;
mem[3805] = 6'b111111;
mem[3806] = 6'b111111;
mem[3807] = 6'b111111;
mem[3808] = 6'b111111;
mem[3809] = 6'b111111;
mem[3810] = 6'b111111;
mem[3811] = 6'b111111;
mem[3812] = 6'b111111;
mem[3813] = 6'b111111;
mem[3814] = 6'b111111;
mem[3815] = 6'b111111;
mem[3816] = 6'b111111;
mem[3817] = 6'b111111;
mem[3818] = 6'b111111;
mem[3819] = 6'b111111;
mem[3820] = 6'b111111;
mem[3821] = 6'b111111;
mem[3822] = 6'b111111;
mem[3823] = 6'b111111;
mem[3824] = 6'b111111;
mem[3825] = 6'b111111;
mem[3826] = 6'b111111;
mem[3827] = 6'b111111;
mem[3828] = 6'b111111;
mem[3829] = 6'b111111;
mem[3830] = 6'b111111;
mem[3831] = 6'b111111;
mem[3832] = 6'b111111;
mem[3833] = 6'b111111;
mem[3834] = 6'b111111;
mem[3835] = 6'b111111;
mem[3836] = 6'b111111;
mem[3837] = 6'b111111;
mem[3838] = 6'b111111;
mem[3839] = 6'b111111;
mem[3840] = 6'b111111;
mem[3841] = 6'b111111;
mem[3842] = 6'b111111;
mem[3843] = 6'b111111;
mem[3844] = 6'b111111;
mem[3845] = 6'b111111;
mem[3846] = 6'b111111;
mem[3847] = 6'b111111;
mem[3848] = 6'b111111;
mem[3849] = 6'b111111;
mem[3850] = 6'b111111;
mem[3851] = 6'b111111;
mem[3852] = 6'b111111;
mem[3853] = 6'b111111;
mem[3854] = 6'b111111;
mem[3855] = 6'b111111;
mem[3856] = 6'b111111;
mem[3857] = 6'b111111;
mem[3858] = 6'b111111;
mem[3859] = 6'b111111;
mem[3860] = 6'b111111;
mem[3861] = 6'b111111;
mem[3862] = 6'b111111;
mem[3863] = 6'b111111;
mem[3864] = 6'b111111;
mem[3865] = 6'b111111;
mem[3866] = 6'b111111;
mem[3867] = 6'b111111;
mem[3868] = 6'b111111;
mem[3869] = 6'b111111;
mem[3870] = 6'b111111;
mem[3871] = 6'b111111;
mem[3872] = 6'b111111;
mem[3873] = 6'b111111;
mem[3874] = 6'b111111;
mem[3875] = 6'b111111;
mem[3876] = 6'b111111;
mem[3877] = 6'b111111;
mem[3878] = 6'b111111;
mem[3879] = 6'b111111;
mem[3880] = 6'b111111;
mem[3881] = 6'b111111;
mem[3882] = 6'b111111;
mem[3883] = 6'b111111;
mem[3884] = 6'b111111;
mem[3885] = 6'b111111;
mem[3886] = 6'b111111;
mem[3887] = 6'b111111;
mem[3888] = 6'b111111;
mem[3889] = 6'b111111;
mem[3890] = 6'b111111;
mem[3891] = 6'b111111;
mem[3892] = 6'b111111;
mem[3893] = 6'b111111;
mem[3894] = 6'b111111;
mem[3895] = 6'b111111;
mem[3896] = 6'b111111;
mem[3897] = 6'b111111;
mem[3898] = 6'b111111;
mem[3899] = 6'b111111;
mem[3900] = 6'b111111;
mem[3901] = 6'b111111;
mem[3902] = 6'b111111;
mem[3903] = 6'b111111;
mem[3904] = 6'b111111;
mem[3905] = 6'b111111;
mem[3906] = 6'b111111;
mem[3907] = 6'b111111;
mem[3908] = 6'b111111;
mem[3909] = 6'b111111;
mem[3910] = 6'b111111;
mem[3911] = 6'b111111;
mem[3912] = 6'b111111;
mem[3913] = 6'b111111;
mem[3914] = 6'b111111;
mem[3915] = 6'b111111;
mem[3916] = 6'b111111;
mem[3917] = 6'b111111;
mem[3918] = 6'b111111;
mem[3919] = 6'b111111;
mem[3920] = 6'b111111;
mem[3921] = 6'b111111;
mem[3922] = 6'b111111;
mem[3923] = 6'b111111;
mem[3924] = 6'b111111;
mem[3925] = 6'b111111;
mem[3926] = 6'b111111;
mem[3927] = 6'b111111;
mem[3928] = 6'b111111;
mem[3929] = 6'b111111;
mem[3930] = 6'b111111;
mem[3931] = 6'b111111;
mem[3932] = 6'b111111;
mem[3933] = 6'b111111;
mem[3934] = 6'b111111;
mem[3935] = 6'b111111;
mem[3936] = 6'b111111;
mem[3937] = 6'b111111;
mem[3938] = 6'b111111;
mem[3939] = 6'b111111;
mem[3940] = 6'b111111;
mem[3941] = 6'b111111;
mem[3942] = 6'b111111;
mem[3943] = 6'b111111;
mem[3944] = 6'b111111;
mem[3945] = 6'b111111;
mem[3946] = 6'b111111;
mem[3947] = 6'b111111;
mem[3948] = 6'b111111;
mem[3949] = 6'b111111;
mem[3950] = 6'b111111;
mem[3951] = 6'b111111;
mem[3952] = 6'b111111;
mem[3953] = 6'b111111;
mem[3954] = 6'b111111;
mem[3955] = 6'b111111;
mem[3956] = 6'b111111;
mem[3957] = 6'b111111;
mem[3958] = 6'b111111;
mem[3959] = 6'b111111;
mem[3960] = 6'b111111;
mem[3961] = 6'b111111;
mem[3962] = 6'b111111;
mem[3963] = 6'b111111;
mem[3964] = 6'b111111;
mem[3965] = 6'b111111;
mem[3966] = 6'b111111;
mem[3967] = 6'b111111;
mem[3968] = 6'b111111;
mem[3969] = 6'b111111;
mem[3970] = 6'b111111;
mem[3971] = 6'b111111;
mem[3972] = 6'b111111;
mem[3973] = 6'b111111;
mem[3974] = 6'b111111;
mem[3975] = 6'b111111;
mem[3976] = 6'b111111;
mem[3977] = 6'b111111;
mem[3978] = 6'b111111;
mem[3979] = 6'b111111;
mem[3980] = 6'b111111;
mem[3981] = 6'b111111;
mem[3982] = 6'b111111;
mem[3983] = 6'b111111;
mem[3984] = 6'b111111;
mem[3985] = 6'b111111;
mem[3986] = 6'b111111;
mem[3987] = 6'b111111;
mem[3988] = 6'b111111;
mem[3989] = 6'b111111;
mem[3990] = 6'b111111;
mem[3991] = 6'b111111;
mem[3992] = 6'b111111;
mem[3993] = 6'b111111;
mem[3994] = 6'b111111;
mem[3995] = 6'b111111;
mem[3996] = 6'b111111;
mem[3997] = 6'b111111;
mem[3998] = 6'b111111;
mem[3999] = 6'b111111;
mem[4000] = 6'b111111;
mem[4001] = 6'b111111;
mem[4002] = 6'b111111;
mem[4003] = 6'b111111;
mem[4004] = 6'b111111;
mem[4005] = 6'b111111;
mem[4006] = 6'b111111;
mem[4007] = 6'b111111;
mem[4008] = 6'b111111;
mem[4009] = 6'b111111;
mem[4010] = 6'b111111;
mem[4011] = 6'b111111;
mem[4012] = 6'b111111;
mem[4013] = 6'b111111;
mem[4014] = 6'b111111;
mem[4015] = 6'b111111;
mem[4016] = 6'b111111;
mem[4017] = 6'b111111;
mem[4018] = 6'b111111;
mem[4019] = 6'b111111;
mem[4020] = 6'b111111;
mem[4021] = 6'b111111;
mem[4022] = 6'b111111;
mem[4023] = 6'b111111;
mem[4024] = 6'b111111;
mem[4025] = 6'b111111;
mem[4026] = 6'b111111;
mem[4027] = 6'b111111;
mem[4028] = 6'b111111;
mem[4029] = 6'b111111;
mem[4030] = 6'b111111;
mem[4031] = 6'b111111;
mem[4032] = 6'b111111;
mem[4033] = 6'b111111;
mem[4034] = 6'b111111;
mem[4035] = 6'b111111;
mem[4036] = 6'b111111;
mem[4037] = 6'b111111;
mem[4038] = 6'b111111;
mem[4039] = 6'b111111;
mem[4040] = 6'b111111;
mem[4041] = 6'b111111;
mem[4042] = 6'b111111;
mem[4043] = 6'b111111;
mem[4044] = 6'b111111;
mem[4045] = 6'b111111;
mem[4046] = 6'b111111;
mem[4047] = 6'b111111;
mem[4048] = 6'b111111;
mem[4049] = 6'b111111;
mem[4050] = 6'b111111;
mem[4051] = 6'b111111;
mem[4052] = 6'b111111;
mem[4053] = 6'b111111;
mem[4054] = 6'b111111;
mem[4055] = 6'b111111;
mem[4056] = 6'b111111;
mem[4057] = 6'b111111;
mem[4058] = 6'b111111;
mem[4059] = 6'b111111;
mem[4060] = 6'b111111;
mem[4061] = 6'b111111;
mem[4062] = 6'b111111;
mem[4063] = 6'b111111;
mem[4064] = 6'b111111;
mem[4065] = 6'b111111;
mem[4066] = 6'b111111;
mem[4067] = 6'b111111;
mem[4068] = 6'b111111;
mem[4069] = 6'b111111;
mem[4070] = 6'b111111;
mem[4071] = 6'b111111;
mem[4072] = 6'b111111;
mem[4073] = 6'b111111;
mem[4074] = 6'b111111;
mem[4075] = 6'b111111;
mem[4076] = 6'b111111;
mem[4077] = 6'b111111;
mem[4078] = 6'b111111;
mem[4079] = 6'b111111;
mem[4080] = 6'b111111;
mem[4081] = 6'b111111;
mem[4082] = 6'b111111;
mem[4083] = 6'b111111;
mem[4084] = 6'b111111;
mem[4085] = 6'b111111;
mem[4086] = 6'b111111;
mem[4087] = 6'b111111;
mem[4088] = 6'b111111;
mem[4089] = 6'b111111;
mem[4090] = 6'b111111;
mem[4091] = 6'b111111;
mem[4092] = 6'b111111;
mem[4093] = 6'b111111;
mem[4094] = 6'b111111;
mem[4095] = 6'b111111;

end

  wire [11:0] addr = {y[6:1], x[6:1]};
  assign pixel = mem[addr][x&11];

endmodule


module palette (
    input  wire [2:0] color_index,
    output wire [5:0] rrggbb
);

  reg [5:0] palette[7:0];

  initial begin
    palette[0] = 6'b001011;  // cyan
    palette[1] = 6'b110110;  // pink
    palette[2] = 6'b101101;  // green
    palette[3] = 6'b111000;  // orange
    palette[4] = 6'b110011;  // purple
    palette[5] = 6'b111100;  // yellow
    palette[6] = 6'b110001;  // red
    palette[7] = 6'b111111;  // white
  end

  assign rrggbb = palette[color_index];

endmodule

/*
Video sync generator, used to drive a VGA monitor.
Timing from: https://en.wikipedia.org/wiki/Video_Graphics_Array
To use:
- Wire the hsync and vsync signals to top level outputs
- Add a 3-bit (or more) "rgb" output to the top level
*/

module vga_sync_generator (
    clk,
    reset,
    hsync,
    vsync,
    display_on,
    hpos,
    vpos
);

  input clk;
  input reset;
  output reg hsync, vsync;
  output display_on;
  output reg [9:0] hpos;
  output reg [9:0] vpos;

  // declarations for TV-simulator sync parameters
  // horizontal constants
  parameter H_DISPLAY = 640;  // horizontal display width
  parameter H_BACK = 48;  // horizontal left border (back porch)
  parameter H_FRONT = 16;  // horizontal right border (front porch)
  parameter H_SYNC = 96;  // horizontal sync width
  // vertical constants
  parameter V_DISPLAY = 480;  // vertical display height
  parameter V_TOP = 33;  // vertical top border
  parameter V_BOTTOM = 10;  // vertical bottom border
  parameter V_SYNC = 2;  // vertical sync # lines
  // derived constants
  parameter H_SYNC_START = H_DISPLAY + H_FRONT;
  parameter H_SYNC_END = H_DISPLAY + H_FRONT + H_SYNC - 1;
  parameter H_MAX = H_DISPLAY + H_BACK + H_FRONT + H_SYNC - 1;
  parameter V_SYNC_START = V_DISPLAY + V_BOTTOM;
  parameter V_SYNC_END = V_DISPLAY + V_BOTTOM + V_SYNC - 1;
  parameter V_MAX = V_DISPLAY + V_TOP + V_BOTTOM + V_SYNC - 1;

  wire hmaxxed = (hpos == H_MAX) || reset;  // set when hpos is maximum
  wire vmaxxed = (vpos == V_MAX) || reset;  // set when vpos is maximum

  // horizontal position counter
  always @(posedge clk) begin
    hsync <= (hpos >= H_SYNC_START && hpos <= H_SYNC_END);
    if (hmaxxed) hpos <= 0;
    else hpos <= hpos + 1;
  end

  // vertical position counter
  always @(posedge clk) begin
    vsync <= (vpos >= V_SYNC_START && vpos <= V_SYNC_END);
    if (hmaxxed)
      if (vmaxxed) vpos <= 0;
      else vpos <= vpos + 1;
  end

  // display_on is set when beam is in "safe" visible frame
  assign display_on = (hpos < H_DISPLAY) && (vpos < V_DISPLAY);

endmodule
